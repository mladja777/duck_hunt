
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017
signal mem : ram_t := (

--			***** COLOR PALLETE *****


	
		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00D4BC00", -- R: 0 G: 188 B: 212
		2 =>	x"001E6933", -- R: 51 G: 105 B: 30
		3 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		4 =>	x"004AC38B", -- R: 139 G: 195 B: 74
		5 =>	x"00205E1B", -- R: 27 G: 94 B: 32
		6 =>	x"000C66A6", -- R: 166 G: 102 B: 12
		7 =>	x"00152A38", -- R: 56 G: 42 B: 21
		--8 =>	x"000A0A0A", -- R: 10 G: 10 B: 10
		--9 =>	x"001A1A1A", -- R: 26 G: 26 B: 26
		--10 =>	x"000B0B0B", -- R: 11 G: 11 B: 11
		8 =>	x"00FFFFFF", -- R: 10 G: 10 B: 10
		9 =>	x"00FFFFFF", -- R: 26 G: 26 B: 26
		10 =>	x"00FFFFFF", -- R: 11 G: 11 B: 11
		11 =>	x"0092CD90", -- R: 144 G: 205 B: 146
		12 =>	x"0050AF4C", -- R: 76 G: 175 B: 80
		13 =>	x"0066B963", -- R: 99 G: 185 B: 102
		14 =>	x"002257FF", -- R: 255 G: 87 B: 34
		15 =>	x"000098FF", -- R: 255 G: 152 B: 0
		16 =>	x"00D7BC07", -- R: 7 G: 188 B: 215
		17 =>	x"00000000", -- Unused
		18 =>	x"00000000", -- Unused
		19 =>	x"00000000", -- Unused
		20 =>	x"00000000", -- Unused
		21 =>	x"00000000", -- Unused
		22 =>	x"00000000", -- Unused
		23 =>	x"00000000", -- Unused
		24 =>	x"00000000", -- Unused
		25 =>	x"00000000", -- Unused
		26 =>	x"00000000", -- Unused
		27 =>	x"00000000", -- Unused
		28 =>	x"00000000", -- Unused
		29 =>	x"00000000", -- Unused
		30 =>	x"00000000", -- Unused
		31 =>	x"00000000", -- Unused
		32 =>	x"00000000", -- Unused
		33 =>	x"00000000", -- Unused
		34 =>	x"00000000", -- Unused
		35 =>	x"00000000", -- Unused
		36 =>	x"00000000", -- Unused
		37 =>	x"00000000", -- Unused
		38 =>	x"00000000", -- Unused
		39 =>	x"00000000", -- Unused
		40 =>	x"00000000", -- Unused
		41 =>	x"00000000", -- Unused
		42 =>	x"00000000", -- Unused
		43 =>	x"00000000", -- Unused
		44 =>	x"00000000", -- Unused
		45 =>	x"00000000", -- Unused
		46 =>	x"00000000", -- Unused
		47 =>	x"00000000", -- Unused
		48 =>	x"00000000", -- Unused
		49 =>	x"00000000", -- Unused
		50 =>	x"00000000", -- Unused
		51 =>	x"00000000", -- Unused
		52 =>	x"00000000", -- Unused
		53 =>	x"00000000", -- Unused
		54 =>	x"00000000", -- Unused
		55 =>	x"00000000", -- Unused
		56 =>	x"00000000", -- Unused
		57 =>	x"00000000", -- Unused
		58 =>	x"00000000", -- Unused
		59 =>	x"00000000", -- Unused
		60 =>	x"00000000", -- Unused
		61 =>	x"00000000", -- Unused
		62 =>	x"00000000", -- Unused
		63 =>	x"00000000", -- Unused
		64 =>	x"00000000", -- Unused
		65 =>	x"00000000", -- Unused
		66 =>	x"00000000", -- Unused
		67 =>	x"00000000", -- Unused
		68 =>	x"00000000", -- Unused
		69 =>	x"00000000", -- Unused
		70 =>	x"00000000", -- Unused
		71 =>	x"00000000", -- Unused
		72 =>	x"00000000", -- Unused
		73 =>	x"00000000", -- Unused
		74 =>	x"00000000", -- Unused
		75 =>	x"00000000", -- Unused
		76 =>	x"00000000", -- Unused
		77 =>	x"00000000", -- Unused
		78 =>	x"00000000", -- Unused
		79 =>	x"00000000", -- Unused
		80 =>	x"00000000", -- Unused
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
		


--			***** 16x16 IMAGES *****


		
		
		

		
		255 =>	x"01010101", -- IMG_16x16_bg00
		256 =>	x"01010101",
		257 =>	x"01010101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01010101",
		261 =>	x"01010101",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01010101",
		265 =>	x"01010101",
		266 =>	x"01010101",
		267 =>	x"01010101",
		268 =>	x"01010101",
		269 =>	x"01010101",
		270 =>	x"01010101",
		271 =>	x"01010101",
		272 =>	x"01020101",
		273 =>	x"01010101",
		274 =>	x"02020101",
		275 =>	x"01010101",
		276 =>	x"01020101",
		277 =>	x"01010101",
		278 =>	x"02020201",
		279 =>	x"01010101",
		280 =>	x"02020203",
		281 =>	x"03010101",
		282 =>	x"01020202",
		283 =>	x"01010101",
		284 =>	x"02040203",
		285 =>	x"03030101",
		286 =>	x"01020202",
		287 =>	x"01010101",
		288 =>	x"02040202",
		289 =>	x"03030303",
		290 =>	x"01010204",
		291 =>	x"01010202",
		292 =>	x"04040402",
		293 =>	x"02030303",
		294 =>	x"01010204",
		295 =>	x"04020204",
		296 =>	x"04040404",
		297 =>	x"02020303",
		298 =>	x"01010204",
		299 =>	x"02020404",
		300 =>	x"04040404",
		301 =>	x"04040203",
		302 =>	x"03010204",
		303 =>	x"02040404",
		304 =>	x"04040404",
		305 =>	x"04040402",
		306 =>	x"03010204",
		307 =>	x"04040404",
		308 =>	x"04040404",
		309 =>	x"04040402",
		310 =>	x"04020204",
		311 =>	x"04040404",
		312 =>	x"04040404",
		313 =>	x"04040404",
		314 =>	x"04040404",
		315 =>	x"04040404",
		316 =>	x"04040404",
		317 =>	x"04040404",
		318 =>	x"04040404",
		319 =>	x"01010101", -- IMG_16x16_bg01
		320 =>	x"01010101",
		321 =>	x"01010101",
		322 =>	x"01010101",
		323 =>	x"01010101",
		324 =>	x"01010101",
		325 =>	x"01010101",
		326 =>	x"01010101",
		327 =>	x"01010101",
		328 =>	x"01010101",
		329 =>	x"01010101",
		330 =>	x"01010101",
		331 =>	x"01010101",
		332 =>	x"01010101",
		333 =>	x"01010101",
		334 =>	x"01010101",
		335 =>	x"01010101",
		336 =>	x"01010101",
		337 =>	x"01010101",
		338 =>	x"01020201",
		339 =>	x"03010101",
		340 =>	x"01010101",
		341 =>	x"01010101",
		342 =>	x"02020101",
		343 =>	x"03030101",
		344 =>	x"01010101",
		345 =>	x"01010102",
		346 =>	x"02030101",
		347 =>	x"02030301",
		348 =>	x"01010101",
		349 =>	x"01010204",
		350 =>	x"02030101",
		351 =>	x"02030303",
		352 =>	x"01010101",
		353 =>	x"01020402",
		354 =>	x"02030101",
		355 =>	x"04020303",
		356 =>	x"03010101",
		357 =>	x"01020402",
		358 =>	x"03030101",
		359 =>	x"04040303",
		360 =>	x"03010101",
		361 =>	x"01040404",
		362 =>	x"02030301",
		363 =>	x"04040203",
		364 =>	x"03030402",
		365 =>	x"04040404",
		366 =>	x"02040301",
		367 =>	x"04040202",
		368 =>	x"03030402",
		369 =>	x"04040404",
		370 =>	x"04040101",
		371 =>	x"04040404",
		372 =>	x"04040404",
		373 =>	x"04040404",
		374 =>	x"04040404",
		375 =>	x"04040404",
		376 =>	x"04040404",
		377 =>	x"04040404",
		378 =>	x"04040404",
		379 =>	x"04040404",
		380 =>	x"04040404",
		381 =>	x"04040404",
		382 =>	x"04040404",
		383 =>	x"01010101", -- IMG_16x16_bg02
		384 =>	x"01010101",
		385 =>	x"01010101",
		386 =>	x"01010101",
		387 =>	x"01010101",
		388 =>	x"01010101",
		389 =>	x"01010101",
		390 =>	x"01010101",
		391 =>	x"01010101",
		392 =>	x"01020101",
		393 =>	x"01010101",
		394 =>	x"01010101",
		395 =>	x"01010101",
		396 =>	x"02020101",
		397 =>	x"01010101",
		398 =>	x"01010102",
		399 =>	x"01010101",
		400 =>	x"02020101",
		401 =>	x"01010101",
		402 =>	x"01010102",
		403 =>	x"01010101",
		404 =>	x"02020101",
		405 =>	x"01010101",
		406 =>	x"01010101",
		407 =>	x"01010101",
		408 =>	x"02020201",
		409 =>	x"01010101",
		410 =>	x"01010101",
		411 =>	x"01010101",
		412 =>	x"02040203",
		413 =>	x"01010101",
		414 =>	x"01010102",
		415 =>	x"01010101",
		416 =>	x"02040203",
		417 =>	x"03010101",
		418 =>	x"01010102",
		419 =>	x"01010101",
		420 =>	x"02040203",
		421 =>	x"03010101",
		422 =>	x"01010102",
		423 =>	x"01010102",
		424 =>	x"02040402",
		425 =>	x"03030101",
		426 =>	x"01010102",
		427 =>	x"01040202",
		428 =>	x"04040402",
		429 =>	x"02040303",
		430 =>	x"01010204",
		431 =>	x"01040404",
		432 =>	x"04040404",
		433 =>	x"02020403",
		434 =>	x"01020404",
		435 =>	x"04040404",
		436 =>	x"04040404",
		437 =>	x"04020204",
		438 =>	x"01020404",
		439 =>	x"04040404",
		440 =>	x"04040404",
		441 =>	x"04040404",
		442 =>	x"04040404",
		443 =>	x"04040404",
		444 =>	x"04040404",
		445 =>	x"04040404",
		446 =>	x"04040404",
		447 =>	x"04040404", -- IMG_16x16_bg10
		448 =>	x"04040404",
		449 =>	x"04040404",
		450 =>	x"04040404",
		451 =>	x"04040404",
		452 =>	x"04040404",
		453 =>	x"04040404",
		454 =>	x"04040404",
		455 =>	x"04040404",
		456 =>	x"04040404",
		457 =>	x"04040404",
		458 =>	x"04040404",
		459 =>	x"04040404",
		460 =>	x"04040404",
		461 =>	x"04040404",
		462 =>	x"04040404",
		463 =>	x"04040404",
		464 =>	x"04040404",
		465 =>	x"04040404",
		466 =>	x"04040404",
		467 =>	x"04040404",
		468 =>	x"04040404",
		469 =>	x"04040404",
		470 =>	x"04040404",
		471 =>	x"04040404",
		472 =>	x"04040404",
		473 =>	x"04040404",
		474 =>	x"04040404",
		475 =>	x"04040404",
		476 =>	x"04040404",
		477 =>	x"04040404",
		478 =>	x"04040404",
		479 =>	x"04040404",
		480 =>	x"04040404",
		481 =>	x"04040404",
		482 =>	x"04040404",
		483 =>	x"04040404",
		484 =>	x"04040404",
		485 =>	x"04040404",
		486 =>	x"04040404",
		487 =>	x"04040404",
		488 =>	x"04040404",
		489 =>	x"04040404",
		490 =>	x"04040404",
		491 =>	x"04040404",
		492 =>	x"04040404",
		493 =>	x"04040404",
		494 =>	x"04040404",
		495 =>	x"04040404",
		496 =>	x"04040404",
		497 =>	x"04040404",
		498 =>	x"04040404",
		499 =>	x"04040404",
		500 =>	x"04040404",
		501 =>	x"04040404",
		502 =>	x"04040404",
		503 =>	x"04040404",
		504 =>	x"04040404",
		505 =>	x"04040404",
		506 =>	x"04040404",
		507 =>	x"04040404",
		508 =>	x"04040404",
		509 =>	x"04040404",
		510 =>	x"04040404",
		511 =>	x"04040404", -- IMG_16x16_bg11
		512 =>	x"04040404",
		513 =>	x"04040404",
		514 =>	x"04040404",
		515 =>	x"04040404",
		516 =>	x"04040404",
		517 =>	x"04040404",
		518 =>	x"04040404",
		519 =>	x"04040404",
		520 =>	x"04040404",
		521 =>	x"04040404",
		522 =>	x"04040404",
		523 =>	x"04040404",
		524 =>	x"04040404",
		525 =>	x"04040504",
		526 =>	x"04040404",
		527 =>	x"04040404",
		528 =>	x"04040404",
		529 =>	x"04040505",
		530 =>	x"04040404",
		531 =>	x"04040404",
		532 =>	x"04040404",
		533 =>	x"04040405",
		534 =>	x"04040404",
		535 =>	x"04040404",
		536 =>	x"04040404",
		537 =>	x"04040405",
		538 =>	x"04040404",
		539 =>	x"04040404",
		540 =>	x"04040404",
		541 =>	x"04040405",
		542 =>	x"04040404",
		543 =>	x"04040404",
		544 =>	x"04040404",
		545 =>	x"04040405",
		546 =>	x"04040404",
		547 =>	x"04040404",
		548 =>	x"04040404",
		549 =>	x"04040505",
		550 =>	x"04040404",
		551 =>	x"04040404",
		552 =>	x"04040404",
		553 =>	x"04040505",
		554 =>	x"04040404",
		555 =>	x"04040404",
		556 =>	x"04040404",
		557 =>	x"04050504",
		558 =>	x"04040404",
		559 =>	x"04040404",
		560 =>	x"04040404",
		561 =>	x"05050404",
		562 =>	x"04040404",
		563 =>	x"04040404",
		564 =>	x"04040404",
		565 =>	x"05050404",
		566 =>	x"04040404",
		567 =>	x"04040404",
		568 =>	x"04040405",
		569 =>	x"05050404",
		570 =>	x"04040404",
		571 =>	x"04040404",
		572 =>	x"04040405",
		573 =>	x"05040404",
		574 =>	x"04040404",
		575 =>	x"04040404", -- IMG_16x16_bg12
		576 =>	x"04040404",
		577 =>	x"04040404",
		578 =>	x"04040404",
		579 =>	x"04040404",
		580 =>	x"04040404",
		581 =>	x"04040404",
		582 =>	x"04040404",
		583 =>	x"04040404",
		584 =>	x"04040404",
		585 =>	x"04040404",
		586 =>	x"04040404",
		587 =>	x"04040404",
		588 =>	x"04040404",
		589 =>	x"04040505",
		590 =>	x"04040404",
		591 =>	x"04040404",
		592 =>	x"04040404",
		593 =>	x"04040405",
		594 =>	x"04040404",
		595 =>	x"04040404",
		596 =>	x"04040404",
		597 =>	x"04040405",
		598 =>	x"04040404",
		599 =>	x"04040404",
		600 =>	x"04040404",
		601 =>	x"04040505",
		602 =>	x"04040404",
		603 =>	x"04040404",
		604 =>	x"04040404",
		605 =>	x"04040505",
		606 =>	x"04040404",
		607 =>	x"04040404",
		608 =>	x"04040404",
		609 =>	x"04040505",
		610 =>	x"04040404",
		611 =>	x"04040404",
		612 =>	x"04040404",
		613 =>	x"04040505",
		614 =>	x"05040404",
		615 =>	x"04040404",
		616 =>	x"04040404",
		617 =>	x"04040405",
		618 =>	x"05040404",
		619 =>	x"04040404",
		620 =>	x"04040404",
		621 =>	x"04040405",
		622 =>	x"05050404",
		623 =>	x"04040404",
		624 =>	x"04040404",
		625 =>	x"04040405",
		626 =>	x"05050404",
		627 =>	x"04040404",
		628 =>	x"04040404",
		629 =>	x"04040404",
		630 =>	x"05050504",
		631 =>	x"04040404",
		632 =>	x"04040404",
		633 =>	x"04040404",
		634 =>	x"04050504",
		635 =>	x"04040404",
		636 =>	x"04040404",
		637 =>	x"04040404",
		638 =>	x"04050404",
		639 =>	x"04040404", -- IMG_16x16_bg20
		640 =>	x"04040404",
		641 =>	x"04040404",
		642 =>	x"04040404",
		643 =>	x"04040404",
		644 =>	x"04040404",
		645 =>	x"04040404",
		646 =>	x"04040404",
		647 =>	x"04040404",
		648 =>	x"04040404",
		649 =>	x"04040404",
		650 =>	x"04040404",
		651 =>	x"04040404",
		652 =>	x"04040404",
		653 =>	x"04040404",
		654 =>	x"04040404",
		655 =>	x"04040404",
		656 =>	x"04040404",
		657 =>	x"04040404",
		658 =>	x"04040404",
		659 =>	x"04040404",
		660 =>	x"04040404",
		661 =>	x"04040404",
		662 =>	x"04040404",
		663 =>	x"04040404",
		664 =>	x"04040404",
		665 =>	x"04040404",
		666 =>	x"04040404",
		667 =>	x"04040404",
		668 =>	x"04040404",
		669 =>	x"04040404",
		670 =>	x"04040404",
		671 =>	x"04040404",
		672 =>	x"04040404",
		673 =>	x"04040404",
		674 =>	x"04040404",
		675 =>	x"04040404",
		676 =>	x"04040404",
		677 =>	x"04040404",
		678 =>	x"04040404",
		679 =>	x"04040404",
		680 =>	x"04040404",
		681 =>	x"04040404",
		682 =>	x"04040404",
		683 =>	x"04040404",
		684 =>	x"04040404",
		685 =>	x"04040404",
		686 =>	x"04040404",
		687 =>	x"04040404",
		688 =>	x"04040404",
		689 =>	x"04040404",
		690 =>	x"04040404",
		691 =>	x"04040404",
		692 =>	x"04040404",
		693 =>	x"04040205",
		694 =>	x"04040404",
		695 =>	x"04040404",
		696 =>	x"04040404",
		697 =>	x"04040405",
		698 =>	x"04040404",
		699 =>	x"04040404",
		700 =>	x"04040404",
		701 =>	x"04040205",
		702 =>	x"04040404",
		703 =>	x"04040404", -- IMG_16x16_bg21
		704 =>	x"04040405",
		705 =>	x"05040404",
		706 =>	x"04040404",
		707 =>	x"04040404",
		708 =>	x"04040405",
		709 =>	x"05040404",
		710 =>	x"04040404",
		711 =>	x"04040404",
		712 =>	x"04040405",
		713 =>	x"05040404",
		714 =>	x"04040404",
		715 =>	x"04040404",
		716 =>	x"04040404",
		717 =>	x"05040404",
		718 =>	x"04040404",
		719 =>	x"04040404",
		720 =>	x"04040405",
		721 =>	x"05040404",
		722 =>	x"04040404",
		723 =>	x"04040404",
		724 =>	x"04040405",
		725 =>	x"04040404",
		726 =>	x"04040404",
		727 =>	x"04040404",
		728 =>	x"04040404",
		729 =>	x"04040404",
		730 =>	x"04040404",
		731 =>	x"04040404",
		732 =>	x"04040404",
		733 =>	x"04040404",
		734 =>	x"04040404",
		735 =>	x"04040404",
		736 =>	x"04040404",
		737 =>	x"04040404",
		738 =>	x"04040404",
		739 =>	x"04040404",
		740 =>	x"04040404",
		741 =>	x"04040404",
		742 =>	x"04040404",
		743 =>	x"04040404",
		744 =>	x"04040404",
		745 =>	x"04040404",
		746 =>	x"04040404",
		747 =>	x"04040404",
		748 =>	x"04040404",
		749 =>	x"04040404",
		750 =>	x"04040404",
		751 =>	x"04040404",
		752 =>	x"04040404",
		753 =>	x"04040404",
		754 =>	x"04040404",
		755 =>	x"04040404",
		756 =>	x"04040404",
		757 =>	x"04040404",
		758 =>	x"04040404",
		759 =>	x"04040404",
		760 =>	x"04040404",
		761 =>	x"04040404",
		762 =>	x"04040404",
		763 =>	x"04040404",
		764 =>	x"04040404",
		765 =>	x"04040404",
		766 =>	x"04040404",
		767 =>	x"04040404", -- IMG_16x16_bg22
		768 =>	x"04040404",
		769 =>	x"04040404",
		770 =>	x"04050404",
		771 =>	x"04040404",
		772 =>	x"04040404",
		773 =>	x"04040404",
		774 =>	x"05050404",
		775 =>	x"04040404",
		776 =>	x"04040404",
		777 =>	x"04040404",
		778 =>	x"05050404",
		779 =>	x"04040404",
		780 =>	x"04040404",
		781 =>	x"04040404",
		782 =>	x"04040404",
		783 =>	x"04040404",
		784 =>	x"04040404",
		785 =>	x"04040404",
		786 =>	x"04040404",
		787 =>	x"04040404",
		788 =>	x"04040404",
		789 =>	x"04040404",
		790 =>	x"04040404",
		791 =>	x"04040404",
		792 =>	x"04040404",
		793 =>	x"04040404",
		794 =>	x"04040404",
		795 =>	x"04040404",
		796 =>	x"04040404",
		797 =>	x"04040404",
		798 =>	x"04040404",
		799 =>	x"04040404",
		800 =>	x"04040404",
		801 =>	x"04040404",
		802 =>	x"04040404",
		803 =>	x"04040404",
		804 =>	x"04040404",
		805 =>	x"04040404",
		806 =>	x"04040404",
		807 =>	x"04040404",
		808 =>	x"04040404",
		809 =>	x"04040404",
		810 =>	x"04040404",
		811 =>	x"04040404",
		812 =>	x"04040404",
		813 =>	x"04040404",
		814 =>	x"04040404",
		815 =>	x"04040404",
		816 =>	x"04040404",
		817 =>	x"04040404",
		818 =>	x"04040404",
		819 =>	x"04040404",
		820 =>	x"04040404",
		821 =>	x"04040404",
		822 =>	x"04040404",
		823 =>	x"05050404",
		824 =>	x"04040404",
		825 =>	x"04040404",
		826 =>	x"04040404",
		827 =>	x"04050204",
		828 =>	x"04040404",
		829 =>	x"04040404",
		830 =>	x"04040404",
		831 =>	x"04040404", -- IMG_16x16_bg30
		832 =>	x"04040404",
		833 =>	x"04020504",
		834 =>	x"04040404",
		835 =>	x"04040404",
		836 =>	x"04040404",
		837 =>	x"04040504",
		838 =>	x"04040404",
		839 =>	x"04040404",
		840 =>	x"04040404",
		841 =>	x"04020504",
		842 =>	x"04040404",
		843 =>	x"04040404",
		844 =>	x"04040404",
		845 =>	x"02050504",
		846 =>	x"04040404",
		847 =>	x"04040404",
		848 =>	x"04040404",
		849 =>	x"05020404",
		850 =>	x"04040404",
		851 =>	x"04040404",
		852 =>	x"04040405",
		853 =>	x"05040404",
		854 =>	x"04040404",
		855 =>	x"04040404",
		856 =>	x"04040405",
		857 =>	x"02040404",
		858 =>	x"04040404",
		859 =>	x"04040404",
		860 =>	x"04040405",
		861 =>	x"02040404",
		862 =>	x"04040404",
		863 =>	x"04040404",
		864 =>	x"04040504",
		865 =>	x"04040404",
		866 =>	x"04040404",
		867 =>	x"04040404",
		868 =>	x"04050504",
		869 =>	x"04040404",
		870 =>	x"04040404",
		871 =>	x"04040404",
		872 =>	x"04050204",
		873 =>	x"04040404",
		874 =>	x"04040404",
		875 =>	x"04040404",
		876 =>	x"04050204",
		877 =>	x"04040404",
		878 =>	x"04040404",
		879 =>	x"04040404",
		880 =>	x"05050404",
		881 =>	x"04040404",
		882 =>	x"04040404",
		883 =>	x"04040404",
		884 =>	x"04040404",
		885 =>	x"04040404",
		886 =>	x"04040404",
		887 =>	x"04040404",
		888 =>	x"04040404",
		889 =>	x"04040404",
		890 =>	x"04040404",
		891 =>	x"04040404",
		892 =>	x"04040404",
		893 =>	x"04040404",
		894 =>	x"04040404",
		895 =>	x"04040404", -- IMG_16x16_bg31
		896 =>	x"04040404",
		897 =>	x"04040404",
		898 =>	x"04040404",
		899 =>	x"04040404",
		900 =>	x"04040404",
		901 =>	x"04040404",
		902 =>	x"04040404",
		903 =>	x"04040404",
		904 =>	x"04040404",
		905 =>	x"04040404",
		906 =>	x"04040404",
		907 =>	x"04040404",
		908 =>	x"04040404",
		909 =>	x"04040404",
		910 =>	x"04040404",
		911 =>	x"04040404",
		912 =>	x"04040404",
		913 =>	x"04040404",
		914 =>	x"04040404",
		915 =>	x"04040404",
		916 =>	x"04040404",
		917 =>	x"04040404",
		918 =>	x"04040404",
		919 =>	x"04040404",
		920 =>	x"04040404",
		921 =>	x"04040404",
		922 =>	x"04040404",
		923 =>	x"04040404",
		924 =>	x"04040404",
		925 =>	x"04040404",
		926 =>	x"04040404",
		927 =>	x"04040404",
		928 =>	x"04040404",
		929 =>	x"04040404",
		930 =>	x"04040404",
		931 =>	x"04040404",
		932 =>	x"04040404",
		933 =>	x"04040404",
		934 =>	x"04040404",
		935 =>	x"04040404",
		936 =>	x"04040404",
		937 =>	x"04040404",
		938 =>	x"04040404",
		939 =>	x"04040404",
		940 =>	x"04040404",
		941 =>	x"04040404",
		942 =>	x"04040404",
		943 =>	x"04040404",
		944 =>	x"04040404",
		945 =>	x"04040404",
		946 =>	x"04040404",
		947 =>	x"04040404",
		948 =>	x"04040404",
		949 =>	x"04040404",
		950 =>	x"04040404",
		951 =>	x"04040404",
		952 =>	x"04040404",
		953 =>	x"04040404",
		954 =>	x"04040404",
		955 =>	x"04040404",
		956 =>	x"04040404",
		957 =>	x"04040404",
		958 =>	x"04040404",
		959 =>	x"04050204", -- IMG_16x16_bg32
		960 =>	x"04040404",
		961 =>	x"04040404",
		962 =>	x"04040404",
		963 =>	x"02050204",
		964 =>	x"04040404",
		965 =>	x"04040404",
		966 =>	x"04040404",
		967 =>	x"04050204",
		968 =>	x"04040404",
		969 =>	x"04040404",
		970 =>	x"04040404",
		971 =>	x"04050204",
		972 =>	x"04040404",
		973 =>	x"04040404",
		974 =>	x"04040404",
		975 =>	x"04050204",
		976 =>	x"04040404",
		977 =>	x"04040404",
		978 =>	x"04040404",
		979 =>	x"04050504",
		980 =>	x"04040404",
		981 =>	x"04040404",
		982 =>	x"04040404",
		983 =>	x"04040504",
		984 =>	x"04040404",
		985 =>	x"04040404",
		986 =>	x"04040404",
		987 =>	x"04040505",
		988 =>	x"04040404",
		989 =>	x"04040404",
		990 =>	x"04040404",
		991 =>	x"04040205",
		992 =>	x"04040404",
		993 =>	x"04040404",
		994 =>	x"04040404",
		995 =>	x"04040405",
		996 =>	x"05040404",
		997 =>	x"04040404",
		998 =>	x"04040404",
		999 =>	x"04040404",
		1000 =>	x"05040404",
		1001 =>	x"04040404",
		1002 =>	x"04040404",
		1003 =>	x"04040404",
		1004 =>	x"05050404",
		1005 =>	x"04040404",
		1006 =>	x"04040404",
		1007 =>	x"04040404",
		1008 =>	x"02050404",
		1009 =>	x"04040404",
		1010 =>	x"04040404",
		1011 =>	x"04040404",
		1012 =>	x"04050404",
		1013 =>	x"04040404",
		1014 =>	x"04040404",
		1015 =>	x"04040404",
		1016 =>	x"04050404",
		1017 =>	x"04040404",
		1018 =>	x"04040404",
		1019 =>	x"04040404",
		1020 =>	x"04050404",
		1021 =>	x"04040404",
		1022 =>	x"04040404",
		1023 =>	x"04040404", -- IMG_16x16_bg40
		1024 =>	x"04040404",
		1025 =>	x"04040404",
		1026 =>	x"04040404",
		1027 =>	x"04040404",
		1028 =>	x"04040404",
		1029 =>	x"04040404",
		1030 =>	x"04040404",
		1031 =>	x"04040404",
		1032 =>	x"04040404",
		1033 =>	x"04040404",
		1034 =>	x"04040404",
		1035 =>	x"04040404",
		1036 =>	x"04040404",
		1037 =>	x"04040404",
		1038 =>	x"04040404",
		1039 =>	x"04040404",
		1040 =>	x"04040404",
		1041 =>	x"04040404",
		1042 =>	x"04040404",
		1043 =>	x"04040404",
		1044 =>	x"04040404",
		1045 =>	x"04040404",
		1046 =>	x"04040404",
		1047 =>	x"04040404",
		1048 =>	x"04040404",
		1049 =>	x"04040404",
		1050 =>	x"04040404",
		1051 =>	x"04040404",
		1052 =>	x"04040404",
		1053 =>	x"04040404",
		1054 =>	x"04040404",
		1055 =>	x"04040404",
		1056 =>	x"04040400",
		1057 =>	x"00040404",
		1058 =>	x"04040404",
		1059 =>	x"04040404",
		1060 =>	x"00000000",
		1061 =>	x"00000000",
		1062 =>	x"04040404",
		1063 =>	x"00000000",
		1064 =>	x"00000606",
		1065 =>	x"06060600",
		1066 =>	x"00000000",
		1067 =>	x"06060606",
		1068 =>	x"06060606",
		1069 =>	x"06060606",
		1070 =>	x"06060606",
		1071 =>	x"06060606",
		1072 =>	x"06060606",
		1073 =>	x"06060606",
		1074 =>	x"06060606",
		1075 =>	x"06060606",
		1076 =>	x"06060606",
		1077 =>	x"06060606",
		1078 =>	x"06060606",
		1079 =>	x"06060606",
		1080 =>	x"06060606",
		1081 =>	x"06060606",
		1082 =>	x"06060606",
		1083 =>	x"06060606",
		1084 =>	x"06060606",
		1085 =>	x"06060606",
		1086 =>	x"06060606",
		1087 =>	x"04040404", -- IMG_16x16_bg41
		1088 =>	x"04040404",
		1089 =>	x"04040404",
		1090 =>	x"04040404",
		1091 =>	x"04040404",
		1092 =>	x"04040404",
		1093 =>	x"04040404",
		1094 =>	x"04040404",
		1095 =>	x"04040404",
		1096 =>	x"04040404",
		1097 =>	x"04040404",
		1098 =>	x"04040404",
		1099 =>	x"04040404",
		1100 =>	x"04040404",
		1101 =>	x"04040404",
		1102 =>	x"04040404",
		1103 =>	x"04040404",
		1104 =>	x"04040404",
		1105 =>	x"04040404",
		1106 =>	x"04040404",
		1107 =>	x"04040404",
		1108 =>	x"04040404",
		1109 =>	x"04040404",
		1110 =>	x"04040404",
		1111 =>	x"04040404",
		1112 =>	x"04040404",
		1113 =>	x"04040404",
		1114 =>	x"04040404",
		1115 =>	x"04040404",
		1116 =>	x"04040404",
		1117 =>	x"04040404",
		1118 =>	x"04040404",
		1119 =>	x"04040404",
		1120 =>	x"04040404",
		1121 =>	x"00040404",
		1122 =>	x"04040404",
		1123 =>	x"04040404",
		1124 =>	x"04000000",
		1125 =>	x"00000004",
		1126 =>	x"04040404",
		1127 =>	x"00000000",
		1128 =>	x"00060606",
		1129 =>	x"06060600",
		1130 =>	x"00000000",
		1131 =>	x"06060606",
		1132 =>	x"06060606",
		1133 =>	x"06060606",
		1134 =>	x"06060606",
		1135 =>	x"06060606",
		1136 =>	x"06060606",
		1137 =>	x"06060606",
		1138 =>	x"06060606",
		1139 =>	x"06060606",
		1140 =>	x"06060606",
		1141 =>	x"06060606",
		1142 =>	x"06060606",
		1143 =>	x"06060606",
		1144 =>	x"06060606",
		1145 =>	x"06060606",
		1146 =>	x"06060606",
		1147 =>	x"06060606",
		1148 =>	x"06060606",
		1149 =>	x"06060606",
		1150 =>	x"06060606",
		1151 =>	x"04040404", -- IMG_16x16_bg42
		1152 =>	x"04050404",
		1153 =>	x"04040404",
		1154 =>	x"04040404",
		1155 =>	x"04040404",
		1156 =>	x"04040404",
		1157 =>	x"04040404",
		1158 =>	x"04040404",
		1159 =>	x"04040404",
		1160 =>	x"04040404",
		1161 =>	x"04040404",
		1162 =>	x"04040404",
		1163 =>	x"04040404",
		1164 =>	x"04040404",
		1165 =>	x"04040404",
		1166 =>	x"04040404",
		1167 =>	x"04040404",
		1168 =>	x"04040404",
		1169 =>	x"04040404",
		1170 =>	x"04040404",
		1171 =>	x"04040404",
		1172 =>	x"04040404",
		1173 =>	x"04040404",
		1174 =>	x"04040404",
		1175 =>	x"04040404",
		1176 =>	x"04040404",
		1177 =>	x"04040404",
		1178 =>	x"04040404",
		1179 =>	x"04040404",
		1180 =>	x"04040404",
		1181 =>	x"04040404",
		1182 =>	x"04040404",
		1183 =>	x"04040404",
		1184 =>	x"00000004",
		1185 =>	x"04040404",
		1186 =>	x"04040404",
		1187 =>	x"00000000",
		1188 =>	x"00000000",
		1189 =>	x"00040404",
		1190 =>	x"04040404",
		1191 =>	x"00060606",
		1192 =>	x"06060606",
		1193 =>	x"00000000",
		1194 =>	x"00000000",
		1195 =>	x"06060606",
		1196 =>	x"06060606",
		1197 =>	x"06060606",
		1198 =>	x"06000006",
		1199 =>	x"06060606",
		1200 =>	x"06060606",
		1201 =>	x"06060606",
		1202 =>	x"06060606",
		1203 =>	x"06060606",
		1204 =>	x"06060606",
		1205 =>	x"06060606",
		1206 =>	x"06060606",
		1207 =>	x"06060606",
		1208 =>	x"06060606",
		1209 =>	x"06060606",
		1210 =>	x"06060606",
		1211 =>	x"06060606",
		1212 =>	x"06060606",
		1213 =>	x"06060606",
		1214 =>	x"06060606",
		1215 =>	x"06060606", -- IMG_16x16_bg50
		1216 =>	x"06060606",
		1217 =>	x"06060606",
		1218 =>	x"06060606",
		1219 =>	x"06060606",
		1220 =>	x"06060606",
		1221 =>	x"06060606",
		1222 =>	x"06060606",
		1223 =>	x"06060606",
		1224 =>	x"06060606",
		1225 =>	x"06060606",
		1226 =>	x"06060606",
		1227 =>	x"06060606",
		1228 =>	x"06060606",
		1229 =>	x"06060606",
		1230 =>	x"06060606",
		1231 =>	x"06060606",
		1232 =>	x"06060606",
		1233 =>	x"06060606",
		1234 =>	x"07070606",
		1235 =>	x"06060606",
		1236 =>	x"06060606",
		1237 =>	x"06060606",
		1238 =>	x"06070707",
		1239 =>	x"06060606",
		1240 =>	x"06060606",
		1241 =>	x"06060606",
		1242 =>	x"06060606",
		1243 =>	x"06060606",
		1244 =>	x"06060606",
		1245 =>	x"06060606",
		1246 =>	x"06060606",
		1247 =>	x"06060606",
		1248 =>	x"06060606",
		1249 =>	x"06060606",
		1250 =>	x"06060607",
		1251 =>	x"06060606",
		1252 =>	x"06060606",
		1253 =>	x"06060606",
		1254 =>	x"06060606",
		1255 =>	x"06060606",
		1256 =>	x"06060606",
		1257 =>	x"06060606",
		1258 =>	x"06060606",
		1259 =>	x"06060606",
		1260 =>	x"06060606",
		1261 =>	x"06060606",
		1262 =>	x"06060606",
		1263 =>	x"06060606",
		1264 =>	x"06060606",
		1265 =>	x"06060606",
		1266 =>	x"06060606",
		1267 =>	x"06060606",
		1268 =>	x"06060606",
		1269 =>	x"06060606",
		1270 =>	x"06060606",
		1271 =>	x"06060606",
		1272 =>	x"06060606",
		1273 =>	x"06060606",
		1274 =>	x"06060606",
		1275 =>	x"06060606",
		1276 =>	x"06060606",
		1277 =>	x"06060606",
		1278 =>	x"06060606",
		1279 =>	x"06060606", -- IMG_16x16_bg51
		1280 =>	x"06060606",
		1281 =>	x"06060606",
		1282 =>	x"06060606",
		1283 =>	x"06060606",
		1284 =>	x"06060606",
		1285 =>	x"06060606",
		1286 =>	x"06060606",
		1287 =>	x"06060606",
		1288 =>	x"06060606",
		1289 =>	x"06060606",
		1290 =>	x"06060606",
		1291 =>	x"06060606",
		1292 =>	x"06060606",
		1293 =>	x"06060606",
		1294 =>	x"06060606",
		1295 =>	x"06060606",
		1296 =>	x"06060606",
		1297 =>	x"06060606",
		1298 =>	x"06060606",
		1299 =>	x"06060606",
		1300 =>	x"06060606",
		1301 =>	x"06060606",
		1302 =>	x"06060606",
		1303 =>	x"06060606",
		1304 =>	x"06060606",
		1305 =>	x"06060606",
		1306 =>	x"06060606",
		1307 =>	x"06060606",
		1308 =>	x"06060606",
		1309 =>	x"06060606",
		1310 =>	x"06060606",
		1311 =>	x"06060606",
		1312 =>	x"06060707",
		1313 =>	x"06060606",
		1314 =>	x"06060606",
		1315 =>	x"06060606",
		1316 =>	x"06060706",
		1317 =>	x"06060606",
		1318 =>	x"06060606",
		1319 =>	x"06060606",
		1320 =>	x"06060606",
		1321 =>	x"06060606",
		1322 =>	x"06060606",
		1323 =>	x"06060606",
		1324 =>	x"06060606",
		1325 =>	x"06060606",
		1326 =>	x"06060606",
		1327 =>	x"06060606",
		1328 =>	x"06060606",
		1329 =>	x"06060606",
		1330 =>	x"06060606",
		1331 =>	x"06060606",
		1332 =>	x"06060606",
		1333 =>	x"06060606",
		1334 =>	x"06060606",
		1335 =>	x"06060606",
		1336 =>	x"06060606",
		1337 =>	x"06060606",
		1338 =>	x"06060606",
		1339 =>	x"06060606",
		1340 =>	x"06060606",
		1341 =>	x"06060606",
		1342 =>	x"06060606",
		1343 =>	x"06060606", -- IMG_16x16_bg52
		1344 =>	x"06060606",
		1345 =>	x"06060606",
		1346 =>	x"06060606",
		1347 =>	x"06060606",
		1348 =>	x"06060606",
		1349 =>	x"06060606",
		1350 =>	x"06060606",
		1351 =>	x"06060606",
		1352 =>	x"06060606",
		1353 =>	x"06060606",
		1354 =>	x"06060607",
		1355 =>	x"06060606",
		1356 =>	x"06060606",
		1357 =>	x"06060606",
		1358 =>	x"06060607",
		1359 =>	x"06060606",
		1360 =>	x"06060606",
		1361 =>	x"06060606",
		1362 =>	x"06060606",
		1363 =>	x"06060606",
		1364 =>	x"06060606",
		1365 =>	x"06060606",
		1366 =>	x"06060606",
		1367 =>	x"06060606",
		1368 =>	x"06060606",
		1369 =>	x"06060606",
		1370 =>	x"06060606",
		1371 =>	x"06060606",
		1372 =>	x"06060606",
		1373 =>	x"06060606",
		1374 =>	x"06060606",
		1375 =>	x"06060606",
		1376 =>	x"06060606",
		1377 =>	x"06060606",
		1378 =>	x"06060606",
		1379 =>	x"06060606",
		1380 =>	x"06060606",
		1381 =>	x"06060606",
		1382 =>	x"06060606",
		1383 =>	x"06060606",
		1384 =>	x"06060606",
		1385 =>	x"06060606",
		1386 =>	x"06060606",
		1387 =>	x"06060606",
		1388 =>	x"06060606",
		1389 =>	x"06060606",
		1390 =>	x"06060606",
		1391 =>	x"06060606",
		1392 =>	x"06060606",
		1393 =>	x"06060606",
		1394 =>	x"06060606",
		1395 =>	x"06060606",
		1396 =>	x"06060606",
		1397 =>	x"06060606",
		1398 =>	x"06060606",
		1399 =>	x"06060606",
		1400 =>	x"06060606",
		1401 =>	x"06060606",
		1402 =>	x"06060606",
		1403 =>	x"06060606",
		1404 =>	x"06060606",
		1405 =>	x"06060606",
		1406 =>	x"06060606",
		1407 =>	x"00000000", -- IMG_16x16_cursor
		1408 =>	x"00000000",
		1409 =>	x"00000000",
		1410 =>	x"00000000",
		1411 =>	x"00000000",
		1412 =>	x"00000008",
		1413 =>	x"00000000",
		1414 =>	x"00000000",
		1415 =>	x"00000000",
		1416 =>	x"00080808",
		1417 =>	x"08080000",
		1418 =>	x"00000000",
		1419 =>	x"00000008",
		1420 =>	x"08080808",
		1421 =>	x"08080808",
		1422 =>	x"00000000",
		1423 =>	x"00000808",
		1424 =>	x"08000008",
		1425 =>	x"00000808",
		1426 =>	x"08000000",
		1427 =>	x"00000808",
		1428 =>	x"00000008",
		1429 =>	x"00000008",
		1430 =>	x"08000000",
		1431 =>	x"00080800",
		1432 =>	x"00000008",
		1433 =>	x"00000000",
		1434 =>	x"08080000",
		1435 =>	x"00080800",
		1436 =>	x"00000008",
		1437 =>	x"00000000",
		1438 =>	x"08080000",
		1439 =>	x"08080809",
		1440 =>	x"0A080808",
		1441 =>	x"08080808",
		1442 =>	x"0A080800",
		1443 =>	x"00080800",
		1444 =>	x"00000008",
		1445 =>	x"00000000",
		1446 =>	x"08080000",
		1447 =>	x"00080800",
		1448 =>	x"00000008",
		1449 =>	x"00000000",
		1450 =>	x"08080000",
		1451 =>	x"00000808",
		1452 =>	x"00000008",
		1453 =>	x"00000008",
		1454 =>	x"08000000",
		1455 =>	x"00000808",
		1456 =>	x"08000008",
		1457 =>	x"00000808",
		1458 =>	x"08000000",
		1459 =>	x"00000008",
		1460 =>	x"08080808",
		1461 =>	x"08080808",
		1462 =>	x"00000000",
		1463 =>	x"00000000",
		1464 =>	x"00080808",
		1465 =>	x"08080000",
		1466 =>	x"00000000",
		1467 =>	x"00000000",
		1468 =>	x"00000008",
		1469 =>	x"00000000",
		1470 =>	x"00000000",
		1471 =>	x"00000000", -- IMG_16x16_pl00
		1472 =>	x"00000000",
		1473 =>	x"00000000",
		1474 =>	x"00000000",
		1475 =>	x"00000000",
		1476 =>	x"00000000",
		1477 =>	x"00000000",
		1478 =>	x"00000000",
		1479 =>	x"00000000",
		1480 =>	x"00000000",
		1481 =>	x"000B0000",
		1482 =>	x"00000000",
		1483 =>	x"00000000",
		1484 =>	x"00000000",
		1485 =>	x"0C0D0C00",
		1486 =>	x"00000000",
		1487 =>	x"00000000",
		1488 =>	x"0E0E000C",
		1489 =>	x"0303030C",
		1490 =>	x"0C000000",
		1491 =>	x"00000000",
		1492 =>	x"0E0E0E0C",
		1493 =>	x"0300030C",
		1494 =>	x"0C000000",
		1495 =>	x"00000000",
		1496 =>	x"000E0E0C",
		1497 =>	x"0303030C",
		1498 =>	x"0C000000",
		1499 =>	x"00000000",
		1500 =>	x"00000E0C",
		1501 =>	x"0C030C0C",
		1502 =>	x"0C000000",
		1503 =>	x"00000000",
		1504 =>	x"0000000C",
		1505 =>	x"0C0C0C0C",
		1506 =>	x"0C0C0000",
		1507 =>	x"00000000",
		1508 =>	x"00000000",
		1509 =>	x"0C0C0C0C",
		1510 =>	x"0C0C0C00",
		1511 =>	x"00000000",
		1512 =>	x"00000000",
		1513 =>	x"000C0C0C",
		1514 =>	x"0C0C0C00",
		1515 =>	x"00000000",
		1516 =>	x"00000000",
		1517 =>	x"000C0C00",
		1518 =>	x"00000000",
		1519 =>	x"00000000",
		1520 =>	x"00000000",
		1521 =>	x"00000008",
		1522 =>	x"08080808",
		1523 =>	x"00000000",
		1524 =>	x"00000000",
		1525 =>	x"00000808",
		1526 =>	x"08080808",
		1527 =>	x"00000000",
		1528 =>	x"00000000",
		1529 =>	x"00000808",
		1530 =>	x"08080808",
		1531 =>	x"00000000",
		1532 =>	x"00000808",
		1533 =>	x"08080808",
		1534 =>	x"08080808",
		1535 =>	x"00000000", -- IMG_16x16_pl01
		1536 =>	x"00000000",
		1537 =>	x"00000000",
		1538 =>	x"00000000",
		1539 =>	x"00000000",
		1540 =>	x"00000000",
		1541 =>	x"00000000",
		1542 =>	x"00000000",
		1543 =>	x"00000000",
		1544 =>	x"00000000",
		1545 =>	x"00000000",
		1546 =>	x"00000000",
		1547 =>	x"00000000",
		1548 =>	x"00000000",
		1549 =>	x"00000000",
		1550 =>	x"00000000",
		1551 =>	x"00000000",
		1552 =>	x"00000000",
		1553 =>	x"00000000",
		1554 =>	x"00000000",
		1555 =>	x"00000000",
		1556 =>	x"00000000",
		1557 =>	x"00000000",
		1558 =>	x"00000000",
		1559 =>	x"00000000",
		1560 =>	x"00000000",
		1561 =>	x"00000000",
		1562 =>	x"00000000",
		1563 =>	x"00000000",
		1564 =>	x"00000000",
		1565 =>	x"00000000",
		1566 =>	x"00000000",
		1567 =>	x"00000000",
		1568 =>	x"00000000",
		1569 =>	x"00000000",
		1570 =>	x"00000000",
		1571 =>	x"00000000",
		1572 =>	x"00000000",
		1573 =>	x"00000000",
		1574 =>	x"00000000",
		1575 =>	x"00000000",
		1576 =>	x"00000000",
		1577 =>	x"00000000",
		1578 =>	x"00000000",
		1579 =>	x"00000000",
		1580 =>	x"00000000",
		1581 =>	x"00000000",
		1582 =>	x"00000000",
		1583 =>	x"00000000",
		1584 =>	x"00000008",
		1585 =>	x"08000000",
		1586 =>	x"00000000",
		1587 =>	x"08000000",
		1588 =>	x"08080808",
		1589 =>	x"08080808",
		1590 =>	x"00000000",
		1591 =>	x"08080808",
		1592 =>	x"08080808",
		1593 =>	x"08080808",
		1594 =>	x"00000000",
		1595 =>	x"08080808",
		1596 =>	x"08080808",
		1597 =>	x"08080000",
		1598 =>	x"00000000",
		1599 =>	x"00000000", -- IMG_16x16_pl10
		1600 =>	x"08080808",
		1601 =>	x"08080808",
		1602 =>	x"08080808",
		1603 =>	x"00000008",
		1604 =>	x"08080808",
		1605 =>	x"08080808",
		1606 =>	x"08080808",
		1607 =>	x"00000808",
		1608 =>	x"08080808",
		1609 =>	x"08080808",
		1610 =>	x"08080808",
		1611 =>	x"00080808",
		1612 =>	x"08080808",
		1613 =>	x"08080808",
		1614 =>	x"08080808",
		1615 =>	x"00000808",
		1616 =>	x"08080808",
		1617 =>	x"08080808",
		1618 =>	x"08080808",
		1619 =>	x"00000008",
		1620 =>	x"08000808",
		1621 =>	x"00080808",
		1622 =>	x"08080808",
		1623 =>	x"00000000",
		1624 =>	x"00000000",
		1625 =>	x"00000000",
		1626 =>	x"08080808",
		1627 =>	x"00000000",
		1628 =>	x"00000000",
		1629 =>	x"00000000",
		1630 =>	x"00080808",
		1631 =>	x"00000000",
		1632 =>	x"00000000",
		1633 =>	x"00000000",
		1634 =>	x"00000808",
		1635 =>	x"00000000",
		1636 =>	x"00000000",
		1637 =>	x"00000000",
		1638 =>	x"00000000",
		1639 =>	x"00000000",
		1640 =>	x"00000000",
		1641 =>	x"00000000",
		1642 =>	x"00000000",
		1643 =>	x"00000000",
		1644 =>	x"00000000",
		1645 =>	x"00000000",
		1646 =>	x"00000000",
		1647 =>	x"00000000",
		1648 =>	x"00000000",
		1649 =>	x"00000000",
		1650 =>	x"00000000",
		1651 =>	x"00000000",
		1652 =>	x"00000000",
		1653 =>	x"00000000",
		1654 =>	x"00000000",
		1655 =>	x"00000000",
		1656 =>	x"00000000",
		1657 =>	x"00000000",
		1658 =>	x"00000000",
		1659 =>	x"00000000",
		1660 =>	x"00000000",
		1661 =>	x"00000000",
		1662 =>	x"00000000",
		1663 =>	x"08080808", -- IMG_16x16_pl11
		1664 =>	x"08080808",
		1665 =>	x"08080000",
		1666 =>	x"00000000",
		1667 =>	x"08080808",
		1668 =>	x"08080808",
		1669 =>	x"08000000",
		1670 =>	x"00000000",
		1671 =>	x"08080808",
		1672 =>	x"08080808",
		1673 =>	x"08000000",
		1674 =>	x"00000000",
		1675 =>	x"08080808",
		1676 =>	x"08080808",
		1677 =>	x"08000000",
		1678 =>	x"00000000",
		1679 =>	x"08080808",
		1680 =>	x"08080808",
		1681 =>	x"08080000",
		1682 =>	x"00000000",
		1683 =>	x"08080808",
		1684 =>	x"08080808",
		1685 =>	x"08080800",
		1686 =>	x"00000000",
		1687 =>	x"08080808",
		1688 =>	x"08080808",
		1689 =>	x"08080800",
		1690 =>	x"00000000",
		1691 =>	x"08080808",
		1692 =>	x"08080808",
		1693 =>	x"08080800",
		1694 =>	x"00000000",
		1695 =>	x"08080808",
		1696 =>	x"08080808",
		1697 =>	x"08000000",
		1698 =>	x"00000000",
		1699 =>	x"00000808",
		1700 =>	x"08000000",
		1701 =>	x"00000000",
		1702 =>	x"00000000",
		1703 =>	x"00000000",
		1704 =>	x"00000000",
		1705 =>	x"00000000",
		1706 =>	x"00000000",
		1707 =>	x"00000000",
		1708 =>	x"0000000E",
		1709 =>	x"0E000000",
		1710 =>	x"00000000",
		1711 =>	x"0000000E",
		1712 =>	x"0E00000E",
		1713 =>	x"0E0E0000",
		1714 =>	x"00000000",
		1715 =>	x"0000000E",
		1716 =>	x"0E0E0000",
		1717 =>	x"0E000000",
		1718 =>	x"00000000",
		1719 =>	x"00000000",
		1720 =>	x"0E0E0E00",
		1721 =>	x"00000000",
		1722 =>	x"00000000",
		1723 =>	x"00000000",
		1724 =>	x"000E0000",
		1725 =>	x"00000000",
		1726 =>	x"00000000",
		1727 =>	x"00000000", -- IMG_16x16_pr00
		1728 =>	x"00000000",
		1729 =>	x"00000000",
		1730 =>	x"00000000",
		1731 =>	x"00000000",
		1732 =>	x"00000000",
		1733 =>	x"00000000",
		1734 =>	x"00000000",
		1735 =>	x"00000000",
		1736 =>	x"00000000",
		1737 =>	x"00000000",
		1738 =>	x"0000000C",
		1739 =>	x"00000000",
		1740 =>	x"00000000",
		1741 =>	x"00000000",
		1742 =>	x"00000C0C",
		1743 =>	x"00000000",
		1744 =>	x"00000000",
		1745 =>	x"00000000",
		1746 =>	x"000C0C0C",
		1747 =>	x"00000000",
		1748 =>	x"00000000",
		1749 =>	x"00000000",
		1750 =>	x"000C0C0C",
		1751 =>	x"00000000",
		1752 =>	x"00000000",
		1753 =>	x"00000000",
		1754 =>	x"000C0C0C",
		1755 =>	x"00000000",
		1756 =>	x"00000000",
		1757 =>	x"00000000",
		1758 =>	x"0C0C0C0C",
		1759 =>	x"00000000",
		1760 =>	x"00000000",
		1761 =>	x"00000000",
		1762 =>	x"0C0C0C0C",
		1763 =>	x"00000000",
		1764 =>	x"00000000",
		1765 =>	x"00000000",
		1766 =>	x"000C0C0C",
		1767 =>	x"00000000",
		1768 =>	x"00000000",
		1769 =>	x"00000000",
		1770 =>	x"000C0C0C",
		1771 =>	x"00000000",
		1772 =>	x"00000000",
		1773 =>	x"00000000",
		1774 =>	x"00000000",
		1775 =>	x"00000000",
		1776 =>	x"00000000",
		1777 =>	x"00000000",
		1778 =>	x"00080808",
		1779 =>	x"00000000",
		1780 =>	x"00080808",
		1781 =>	x"00000000",
		1782 =>	x"08080808",
		1783 =>	x"00080808",
		1784 =>	x"08080808",
		1785 =>	x"08080808",
		1786 =>	x"08080808",
		1787 =>	x"00000808",
		1788 =>	x"08080808",
		1789 =>	x"08080808",
		1790 =>	x"08080808",
		1791 =>	x"00000000", -- IMG_16x16_pr01
		1792 =>	x"00000000",
		1793 =>	x"00000000",
		1794 =>	x"00000000",
		1795 =>	x"00000000",
		1796 =>	x"00000000",
		1797 =>	x"00000000",
		1798 =>	x"00000000",
		1799 =>	x"0C0C0000",
		1800 =>	x"00000000",
		1801 =>	x"00000000",
		1802 =>	x"00000000",
		1803 =>	x"0C030C0C",
		1804 =>	x"00000F0F",
		1805 =>	x"00000000",
		1806 =>	x"00000000",
		1807 =>	x"0303030C",
		1808 =>	x"0C0F0F0F",
		1809 =>	x"00000000",
		1810 =>	x"00000000",
		1811 =>	x"0300030C",
		1812 =>	x"0C0F0F0F",
		1813 =>	x"00000000",
		1814 =>	x"00000000",
		1815 =>	x"0303030C",
		1816 =>	x"0C0F0F00",
		1817 =>	x"00000000",
		1818 =>	x"00000000",
		1819 =>	x"0C030C0C",
		1820 =>	x"0C0F0000",
		1821 =>	x"00000000",
		1822 =>	x"00000000",
		1823 =>	x"0C0C0C0C",
		1824 =>	x"0C000000",
		1825 =>	x"00000000",
		1826 =>	x"00000000",
		1827 =>	x"0C0C0C0C",
		1828 =>	x"0C000000",
		1829 =>	x"00000000",
		1830 =>	x"00000000",
		1831 =>	x"0C0C0C0C",
		1832 =>	x"00000000",
		1833 =>	x"00000000",
		1834 =>	x"00000000",
		1835 =>	x"00000C00",
		1836 =>	x"00000000",
		1837 =>	x"00000000",
		1838 =>	x"00000000",
		1839 =>	x"08000000",
		1840 =>	x"00000000",
		1841 =>	x"00000000",
		1842 =>	x"00000000",
		1843 =>	x"08080800",
		1844 =>	x"00000000",
		1845 =>	x"00000000",
		1846 =>	x"00000000",
		1847 =>	x"08080808",
		1848 =>	x"00000000",
		1849 =>	x"00000000",
		1850 =>	x"00000000",
		1851 =>	x"08080808",
		1852 =>	x"08080808",
		1853 =>	x"00000000",
		1854 =>	x"00000000",
		1855 =>	x"00000808", -- IMG_16x16_pr10
		1856 =>	x"08080808",
		1857 =>	x"08080808",
		1858 =>	x"08080808",
		1859 =>	x"00000008",
		1860 =>	x"08080808",
		1861 =>	x"08080808",
		1862 =>	x"08080808",
		1863 =>	x"00000008",
		1864 =>	x"08080808",
		1865 =>	x"08080808",
		1866 =>	x"08080808",
		1867 =>	x"00000000",
		1868 =>	x"00080808",
		1869 =>	x"08080808",
		1870 =>	x"08080808",
		1871 =>	x"00000000",
		1872 =>	x"00000808",
		1873 =>	x"08080808",
		1874 =>	x"08080808",
		1875 =>	x"00000000",
		1876 =>	x"00000008",
		1877 =>	x"08080808",
		1878 =>	x"08080808",
		1879 =>	x"00000000",
		1880 =>	x"00000008",
		1881 =>	x"08080808",
		1882 =>	x"08080808",
		1883 =>	x"00000000",
		1884 =>	x"00000808",
		1885 =>	x"08080808",
		1886 =>	x"08080808",
		1887 =>	x"00000000",
		1888 =>	x"00000808",
		1889 =>	x"08080808",
		1890 =>	x"08080800",
		1891 =>	x"00000000",
		1892 =>	x"00080808",
		1893 =>	x"08080808",
		1894 =>	x"00000000",
		1895 =>	x"00000000",
		1896 =>	x"00000808",
		1897 =>	x"08080000",
		1898 =>	x"00000000",
		1899 =>	x"00000000",
		1900 =>	x"00000000",
		1901 =>	x"0000000E",
		1902 =>	x"0E000000",
		1903 =>	x"00000000",
		1904 =>	x"0000000E",
		1905 =>	x"0E000E0E",
		1906 =>	x"0E000000",
		1907 =>	x"00000000",
		1908 =>	x"00000E0E",
		1909 =>	x"0E000E0E",
		1910 =>	x"0E000000",
		1911 =>	x"00000000",
		1912 =>	x"0000000E",
		1913 =>	x"0000000E",
		1914 =>	x"00000000",
		1915 =>	x"00000000",
		1916 =>	x"00000000",
		1917 =>	x"00000000",
		1918 =>	x"00000000",
		1919 =>	x"08080808", -- IMG_16x16_pr11
		1920 =>	x"08080808",
		1921 =>	x"08080000",
		1922 =>	x"00000000",
		1923 =>	x"08080808",
		1924 =>	x"08080808",
		1925 =>	x"08080800",
		1926 =>	x"00000000",
		1927 =>	x"08080808",
		1928 =>	x"08080808",
		1929 =>	x"08080808",
		1930 =>	x"08000000",
		1931 =>	x"08080808",
		1932 =>	x"08080808",
		1933 =>	x"08080808",
		1934 =>	x"08080000",
		1935 =>	x"08080808",
		1936 =>	x"08080808",
		1937 =>	x"08080808",
		1938 =>	x"08080800",
		1939 =>	x"08080808",
		1940 =>	x"08080808",
		1941 =>	x"08080808",
		1942 =>	x"00000000",
		1943 =>	x"08080800",
		1944 =>	x"00080808",
		1945 =>	x"08080000",
		1946 =>	x"00000000",
		1947 =>	x"08000000",
		1948 =>	x"00000008",
		1949 =>	x"00000000",
		1950 =>	x"00000000",
		1951 =>	x"00000000",
		1952 =>	x"00000000",
		1953 =>	x"00000000",
		1954 =>	x"00000000",
		1955 =>	x"00000000",
		1956 =>	x"00000000",
		1957 =>	x"00000000",
		1958 =>	x"00000000",
		1959 =>	x"00000000",
		1960 =>	x"00000000",
		1961 =>	x"00000000",
		1962 =>	x"00000000",
		1963 =>	x"00000000",
		1964 =>	x"00000000",
		1965 =>	x"00000000",
		1966 =>	x"00000000",
		1967 =>	x"00000000",
		1968 =>	x"00000000",
		1969 =>	x"00000000",
		1970 =>	x"00000000",
		1971 =>	x"00000000",
		1972 =>	x"00000000",
		1973 =>	x"00000000",
		1974 =>	x"00000000",
		1975 =>	x"00000000",
		1976 =>	x"00000000",
		1977 =>	x"00000000",
		1978 =>	x"00000000",
		1979 =>	x"00000000",
		1980 =>	x"00000000",
		1981 =>	x"00000000",
		1982 =>	x"00000000",
		1983 =>	x"10010101", -- IMG_16x16_sky
		1984 =>	x"01010101",
		1985 =>	x"01010101",
		1986 =>	x"01010101",
		1987 =>	x"01010101",
		1988 =>	x"01010101",
		1989 =>	x"01010101",
		1990 =>	x"01010101",
		1991 =>	x"01010101",
		1992 =>	x"01010101",
		1993 =>	x"01010101",
		1994 =>	x"01010101",
		1995 =>	x"01010101",
		1996 =>	x"01010101",
		1997 =>	x"01010101",
		1998 =>	x"01010101",
		1999 =>	x"01010101",
		2000 =>	x"01010101",
		2001 =>	x"01010101",
		2002 =>	x"01010101",
		2003 =>	x"01010101",
		2004 =>	x"01010101",
		2005 =>	x"01010101",
		2006 =>	x"01010101",
		2007 =>	x"01010101",
		2008 =>	x"01010101",
		2009 =>	x"01010101",
		2010 =>	x"01010101",
		2011 =>	x"01010101",
		2012 =>	x"01010101",
		2013 =>	x"01010101",
		2014 =>	x"01010101",
		2015 =>	x"01010101",
		2016 =>	x"01010101",
		2017 =>	x"01010101",
		2018 =>	x"01010101",
		2019 =>	x"01010101",
		2020 =>	x"01010101",
		2021 =>	x"01010101",
		2022 =>	x"01010101",
		2023 =>	x"01010101",
		2024 =>	x"01010101",
		2025 =>	x"01010101",
		2026 =>	x"01010101",
		2027 =>	x"01010101",
		2028 =>	x"01010101",
		2029 =>	x"01010101",
		2030 =>	x"01010101",
		2031 =>	x"01010101",
		2032 =>	x"01010101",
		2033 =>	x"01010101",
		2034 =>	x"01010101",
		2035 =>	x"01010101",
		2036 =>	x"01010101",
		2037 =>	x"01010101",
		2038 =>	x"01010101",
		2039 =>	x"01010101",
		2040 =>	x"01010101",
		2041 =>	x"01010101",
		2042 =>	x"01010101",
		2043 =>	x"01010101",
		2044 =>	x"01010101",
		2045 =>	x"01010101",
		2046 =>	x"01010101",
--			***** MAP *****

		2047 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2048 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2049 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2050 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2051 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2052 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2053 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2054 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2055 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2056 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2057 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2058 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2059 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2060 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2061 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2062 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2063 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2064 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2065 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2066 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2067 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2068 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2069 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2070 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2071 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2072 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2073 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2074 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2075 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2076 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2077 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2078 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2079 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2080 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2081 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2082 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2083 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2084 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2085 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2086 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2087 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2088 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2089 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2090 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2091 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2092 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2093 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2094 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2095 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2096 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2097 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2098 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2099 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2100 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2101 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2102 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2103 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2104 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2105 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2106 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2107 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2108 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2109 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2110 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2111 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2112 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2113 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2114 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2115 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2116 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2117 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2118 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2119 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2120 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2121 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2122 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2123 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2124 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2125 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2126 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2127 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2128 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2129 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2130 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2131 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2132 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2133 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2134 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2135 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2136 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2137 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2138 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2139 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2140 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2141 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2142 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2143 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2144 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2145 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2146 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2147 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2148 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2149 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2150 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2151 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2152 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2153 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2154 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2155 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2156 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2157 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2158 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2159 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2160 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2161 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2162 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2163 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2164 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2165 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2166 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2167 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2168 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2169 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2170 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2171 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2172 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2173 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2174 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2175 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2176 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2177 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2178 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2179 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2180 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2181 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2182 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2183 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2184 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2185 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2186 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2187 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2188 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2189 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2190 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2191 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2192 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2193 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2194 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2195 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2196 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2197 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2198 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2199 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2200 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2201 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2202 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2203 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2204 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2205 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2206 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2207 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2208 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2209 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2210 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2211 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2212 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2213 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2214 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2215 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2216 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2217 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2218 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2219 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2220 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2221 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2222 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2223 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2224 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2225 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2226 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2227 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2228 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2229 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2230 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2231 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2232 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2233 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2234 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2235 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2236 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2237 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2238 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2239 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2240 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2241 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2242 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2243 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2244 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2245 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2246 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2247 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2248 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2249 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2250 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2251 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2252 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2253 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2254 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2255 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2256 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2257 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2258 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2259 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2260 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2261 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2262 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2263 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2264 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2265 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2266 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2267 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2268 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2269 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2270 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2271 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2272 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2273 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2274 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2275 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2276 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2277 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2278 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2279 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2280 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2281 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2282 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2283 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2284 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2285 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2286 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2287 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2288 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2289 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2290 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2291 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2292 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2293 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2294 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2295 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2296 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2297 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2298 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2299 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2300 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2301 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2302 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2303 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2304 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2305 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2306 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2307 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2308 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2309 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2310 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2311 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2312 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2313 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2314 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2315 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2316 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2317 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2318 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2319 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2320 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2321 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2322 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2323 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2324 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2325 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2326 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2327 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2328 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2329 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2330 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2331 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2332 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2333 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2334 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2335 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2336 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2337 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2338 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2339 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2340 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2341 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2342 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2343 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2344 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2345 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2346 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2347 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2348 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2349 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2350 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2351 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2352 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2353 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2354 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2355 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2356 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2357 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2358 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2359 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2360 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2361 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2362 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2363 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2364 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2365 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2366 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2367 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2368 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2369 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2370 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2371 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2372 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2373 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2374 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2375 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2376 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2377 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2378 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2379 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2380 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2381 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2382 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2383 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2384 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2385 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2386 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2387 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2388 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2389 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2390 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2391 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2392 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2393 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2394 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2395 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2396 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2397 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2398 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2399 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2400 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2401 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2402 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2403 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2404 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2405 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2406 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2407 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2408 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2409 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2410 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2411 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2412 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2413 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2414 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2415 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2416 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2417 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2418 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2419 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2420 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2421 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2422 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2423 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2424 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2425 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2426 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2427 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2428 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2429 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2430 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2431 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2432 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2433 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2434 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2435 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2436 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2437 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2438 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2439 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2440 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2441 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2442 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2443 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2444 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2445 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2446 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2447 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2448 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2449 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2450 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2451 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2452 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2453 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2454 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2455 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2456 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2457 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2458 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2459 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2460 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2461 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2462 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2463 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2464 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2465 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2466 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2467 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2468 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2469 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2470 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2471 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2472 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2473 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2474 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2475 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2476 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2477 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2478 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2479 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2480 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2481 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2482 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2483 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2484 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2485 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2486 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2487 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2488 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2489 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2490 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2491 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2492 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2493 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2494 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2495 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2496 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2497 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2498 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2499 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2500 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2501 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2502 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2503 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2504 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2505 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2506 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2507 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2508 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2509 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2510 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2511 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2512 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2513 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2514 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2515 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2516 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2517 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2518 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2519 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2520 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2521 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2522 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2523 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2524 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2525 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2526 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2527 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2528 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2529 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2530 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2531 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2532 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2533 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2534 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2535 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2536 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2537 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2538 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2539 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2540 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2541 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2542 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2543 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2544 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2545 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2546 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2547 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2548 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2549 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2550 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2551 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2552 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2553 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2554 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2555 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2556 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2557 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2558 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2559 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2560 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2561 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2562 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2563 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2564 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2565 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2566 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2567 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2568 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2569 =>	x"000007BF", -- z: 0 rsot: 0 ptr: 1983
		2570 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2571 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2572 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2573 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2574 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2575 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2576 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2577 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2578 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2579 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2580 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2581 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2582 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2583 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2584 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2585 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2586 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2587 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2588 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2589 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2590 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2591 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2592 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2593 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2594 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2595 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2596 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2597 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2598 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2599 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2600 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2601 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2602 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2603 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2604 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2605 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2606 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2607 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2608 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2609 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2610 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2611 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2612 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2613 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2614 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2615 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2616 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2617 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2618 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2619 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2620 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2621 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2622 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2623 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2624 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2625 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2626 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2627 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2628 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2629 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2630 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2631 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2632 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2633 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2634 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2635 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2636 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2637 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2638 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2639 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2640 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2641 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2642 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2643 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2644 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2645 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2646 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2647 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2648 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2649 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2650 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2651 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2652 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2653 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2654 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2655 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2656 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2657 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2658 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2659 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2660 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2661 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2662 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2663 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2664 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2665 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2666 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2667 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2668 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2669 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2670 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2671 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2672 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2673 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2674 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2675 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2676 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2677 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2678 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2679 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2680 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2681 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2682 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2683 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2684 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2685 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2686 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2687 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2688 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2689 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2690 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2691 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2692 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2693 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2694 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2695 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2696 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2697 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2698 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2699 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2700 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2701 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2702 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2703 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2704 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2705 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2706 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2707 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2708 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2709 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2710 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2711 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2712 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2713 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2714 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2715 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2716 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2717 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2718 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2719 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2720 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2721 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2722 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2723 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2724 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2725 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2726 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2727 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2728 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2729 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2730 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2731 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2732 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2733 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2734 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2735 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2736 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2737 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2738 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2739 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2740 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2741 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2742 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2743 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2744 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2745 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2746 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2747 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2748 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2749 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2750 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2751 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2752 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2753 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2754 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2755 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2756 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2757 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2758 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2759 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2760 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2761 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2762 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2763 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2764 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2765 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2766 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2767 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2768 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2769 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2770 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2771 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2772 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2773 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2774 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2775 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2776 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2777 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2778 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2779 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2780 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2781 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2782 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2783 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2784 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2785 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2786 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2787 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2788 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2789 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2790 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2791 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2792 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2793 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2794 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2795 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2796 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2797 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2798 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2799 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2800 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2801 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2802 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2803 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2804 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2805 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2806 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2807 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2808 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2809 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2810 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2811 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2812 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2813 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2814 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2815 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2816 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2817 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2818 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2819 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2820 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2821 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2822 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2823 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2824 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2825 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2826 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2827 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2828 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2829 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2830 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2831 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2832 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2833 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2834 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2835 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2836 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2837 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2838 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2839 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2840 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2841 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2842 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2843 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2844 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2845 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2846 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2847 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2848 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2849 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2850 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2851 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2852 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2853 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2854 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2855 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2856 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2857 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2858 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2859 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2860 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2861 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2862 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2863 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2864 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2865 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2866 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2867 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2868 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2869 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2870 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2871 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2872 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2873 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2874 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2875 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2876 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2877 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2878 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2879 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2880 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2881 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2882 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2883 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2884 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2885 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2886 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2887 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2888 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2889 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2890 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2891 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2892 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2893 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2894 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2895 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2896 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2897 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2898 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2899 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2900 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2901 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2902 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2903 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2904 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2905 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2906 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2907 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2908 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2909 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2910 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2911 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2912 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2913 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2914 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2915 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2916 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2917 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2918 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2919 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2920 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2921 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2922 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2923 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2924 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2925 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2926 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2927 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2928 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2929 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2930 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2931 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2932 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2933 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2934 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2935 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2936 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2937 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2938 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2939 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2940 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2941 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2942 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2943 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2944 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2945 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2946 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2947 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2948 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2949 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2950 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2951 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2952 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2953 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2954 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2955 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2956 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2957 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2958 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2959 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2960 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2961 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2962 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2963 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2964 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2965 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2966 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2967 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2968 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2969 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2970 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2971 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2972 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2973 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2974 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2975 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2976 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2977 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2978 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2979 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2980 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2981 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2982 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2983 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2984 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2985 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2986 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2987 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2988 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2989 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2990 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2991 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2992 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2993 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2994 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2995 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2996 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2997 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2998 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		2999 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3000 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3001 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3002 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3003 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3004 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3005 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3006 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3007 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3008 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3009 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3010 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3011 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3012 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3013 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3014 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3015 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3016 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3017 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3018 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3019 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3020 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3021 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3022 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3023 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3024 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3025 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3026 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3027 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3028 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3029 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3030 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3031 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3032 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3033 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3034 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3035 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3036 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3037 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3038 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3039 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3040 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3041 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3042 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3043 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3044 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3045 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3046 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3047 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3048 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3049 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3050 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3051 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3052 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3053 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3054 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3055 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3056 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3057 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3058 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3059 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3060 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3061 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3062 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3063 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3064 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3065 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3066 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3067 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3068 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3069 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3070 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3071 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3072 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3073 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3074 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3075 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3076 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3077 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3078 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3079 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3080 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3081 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3082 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3083 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3084 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3085 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3086 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3087 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3088 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3089 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3090 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3091 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3092 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3093 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3094 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3095 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3096 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3097 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3098 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3099 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3100 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3101 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3102 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3103 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3104 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3105 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3106 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3107 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3108 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3109 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3110 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3111 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3112 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3113 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3114 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3115 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3116 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3117 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3118 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3119 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3120 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3121 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3122 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3123 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3124 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3125 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3126 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3127 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3128 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3129 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3130 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3131 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3132 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3133 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3134 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3135 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3136 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3137 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3138 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3139 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3140 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3141 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3142 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3143 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3144 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3145 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3146 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3147 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3148 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3149 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3150 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3151 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3152 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3153 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3154 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3155 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3156 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3157 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3158 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3159 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3160 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3161 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3162 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3163 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3164 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3165 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3166 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3167 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3168 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3169 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3170 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3171 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3172 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3173 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3174 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3175 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3176 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3177 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3178 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3179 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3180 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3181 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3182 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3183 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3184 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3185 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3186 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3187 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3188 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3189 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3190 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3191 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3192 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3193 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3194 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3195 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3196 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3197 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3198 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3199 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3200 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3201 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3202 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3203 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3204 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3205 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3206 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3207 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3208 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3209 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3210 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3211 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3212 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3213 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3214 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3215 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3216 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3217 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3218 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3219 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3220 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3221 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3222 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3223 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3224 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3225 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3226 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3227 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3228 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3229 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3230 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3231 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3232 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3233 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3234 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3235 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3236 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3237 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3238 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3239 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3240 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3241 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3242 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3243 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3244 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3245 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3246 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3247 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3248 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3249 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3250 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3251 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3252 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3253 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3254 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3255 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3256 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3257 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3258 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3259 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3260 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3261 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3262 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3263 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3264 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3265 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3266 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3267 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3268 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3269 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3270 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3271 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3272 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3273 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3274 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3275 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3276 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3277 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3278 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3279 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3280 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3281 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3282 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3283 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3284 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3285 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3286 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3287 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3288 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3289 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3290 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3291 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3292 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3293 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3294 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3295 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3296 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3297 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3298 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3299 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3300 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3301 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3302 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3303 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3304 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3305 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3306 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3307 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3308 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3309 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3310 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3311 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3312 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3313 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3314 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3315 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3316 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3317 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3318 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3319 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3320 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3321 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3322 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3323 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3324 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3325 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3326 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3327 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3328 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3329 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3330 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3331 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3332 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3333 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3334 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3335 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3336 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3337 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3338 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3339 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3340 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3341 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3342 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3343 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3344 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3345 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3346 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3347 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3348 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3349 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3350 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3351 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3352 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3353 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3354 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3355 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3356 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3357 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3358 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3359 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3360 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3361 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3362 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3363 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3364 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3365 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3366 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3367 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3368 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3369 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3370 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3371 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3372 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3373 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3374 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3375 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3376 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3377 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3378 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3379 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3380 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3381 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3382 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3383 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3384 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3385 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3386 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3387 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3388 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3389 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3390 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3391 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3392 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3393 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3394 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3395 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3396 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3397 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3398 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3399 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3400 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3401 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3402 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3403 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3404 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3405 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3406 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3407 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3408 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3409 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3410 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3411 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3412 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3413 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3414 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3415 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3416 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3417 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3418 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3419 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3420 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3421 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3422 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3423 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3424 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3425 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3426 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3427 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3428 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3429 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3430 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3431 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3432 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3433 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3434 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3435 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3436 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3437 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3438 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3439 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3440 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3441 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3442 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3443 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3444 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3445 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3446 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3447 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3448 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3449 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3450 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3451 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3452 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3453 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3454 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3455 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3456 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3457 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3458 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3459 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3460 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3461 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3462 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3463 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3464 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3465 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3466 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3467 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3468 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3469 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3470 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3471 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3472 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3473 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3474 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3475 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3476 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3477 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3478 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3479 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3480 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3481 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3482 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3483 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3484 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3485 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3486 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3487 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3488 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3489 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3490 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3491 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3492 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3493 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3494 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3495 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3496 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3497 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3498 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3499 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3500 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3501 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3502 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3503 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3504 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3505 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3506 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3507 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3508 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3509 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3510 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3511 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3512 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3513 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3514 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3515 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3516 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3517 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3518 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3519 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3520 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3521 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3522 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3523 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3524 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3525 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3526 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3527 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3528 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3529 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3530 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3531 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3532 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3533 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3534 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3535 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3536 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3537 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3538 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3539 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3540 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3541 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3542 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3543 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3544 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3545 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3546 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3547 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3548 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3549 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3550 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3551 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3552 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3553 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3554 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3555 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3556 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3557 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3558 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3559 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3560 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3561 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3562 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3563 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3564 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3565 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3566 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3567 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3568 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3569 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3570 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3571 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3572 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3573 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3574 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3575 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3576 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3577 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3578 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3579 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3580 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3581 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3582 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3583 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3584 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3585 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3586 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3587 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3588 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3589 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3590 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3591 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3592 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3593 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3594 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3595 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3596 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3597 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3598 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3599 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3600 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3601 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3602 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3603 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3604 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3605 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3606 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3607 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3608 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3609 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3610 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3611 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3612 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3613 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3614 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3615 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3616 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3617 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3618 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3619 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3620 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3621 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3622 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3623 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3624 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3625 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3626 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3627 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3628 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3629 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3630 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3631 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3632 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3633 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3634 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3635 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3636 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3637 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3638 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3639 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3640 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3641 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3642 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3643 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3644 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3645 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3646 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3647 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3648 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3649 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3650 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3651 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3652 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3653 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3654 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3655 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3656 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3657 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3658 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3659 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3660 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3661 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3662 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3663 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3664 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3665 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3666 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3667 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3668 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3669 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3670 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3671 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3672 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3673 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3674 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3675 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3676 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3677 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3678 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3679 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3680 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3681 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3682 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3683 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3684 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3685 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3686 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3687 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3688 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3689 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3690 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3691 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3692 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3693 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3694 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3695 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3696 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3697 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3698 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3699 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3700 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3701 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3702 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3703 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3704 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3705 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3706 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3707 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3708 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3709 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3710 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3711 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3712 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3713 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3714 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3715 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3716 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3717 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3718 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3719 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3720 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3721 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3722 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3723 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3724 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3725 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3726 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3727 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3728 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3729 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3730 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3731 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3732 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3733 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3734 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3735 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3736 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3737 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3738 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3739 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3740 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3741 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3742 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3743 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3744 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3745 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3746 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3747 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3748 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3749 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3750 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3751 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3752 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3753 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3754 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3755 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3756 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3757 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3758 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3759 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3760 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3761 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3762 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3763 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3764 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3765 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3766 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3767 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3768 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3769 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3770 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3771 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3772 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3773 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3774 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3775 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3776 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3777 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3778 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3779 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3780 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3781 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3782 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3783 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3784 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3785 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3786 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3787 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3788 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3789 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3790 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3791 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3792 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3793 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3794 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3795 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3796 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3797 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3798 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3799 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3800 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3801 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3802 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3803 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3804 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3805 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3806 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3807 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3808 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3809 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3810 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3811 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3812 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3813 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3814 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3815 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3816 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3817 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3818 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3819 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3820 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3821 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3822 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3823 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3824 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3825 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3826 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3827 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3828 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3829 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3830 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3831 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3832 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3833 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3834 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3835 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3836 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3837 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3838 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3839 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3840 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3841 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3842 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3843 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3844 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3845 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3846 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3847 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3848 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3849 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3850 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3851 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3852 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3853 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3854 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3855 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3856 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3857 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3858 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3859 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3860 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3861 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3862 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3863 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3864 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3865 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3866 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3867 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3868 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3869 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3870 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3871 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3872 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3873 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3874 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3875 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3876 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3877 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3878 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3879 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3880 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3881 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3882 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3883 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3884 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3885 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3886 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3887 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3888 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3889 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3890 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3891 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3892 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3893 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3894 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3895 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3896 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3897 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3898 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3899 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3900 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3901 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3902 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3903 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3904 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3905 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3906 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3907 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3908 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3909 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3910 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3911 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3912 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3913 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3914 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3915 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3916 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3917 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3918 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3919 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3920 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3921 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3922 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3923 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3924 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3925 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3926 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3927 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3928 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3929 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3930 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3931 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3932 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3933 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3934 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3935 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3936 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3937 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3938 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3939 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3940 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3941 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3942 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3943 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3944 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3945 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3946 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3947 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3948 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3949 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3950 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3951 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3952 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3953 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3954 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3955 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3956 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3957 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3958 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3959 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3960 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3961 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3962 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3963 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3964 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3965 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3966 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3967 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3968 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3969 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3970 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3971 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3972 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3973 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3974 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3975 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3976 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3977 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3978 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3979 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3980 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3981 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3982 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3983 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3984 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3985 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3986 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3987 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3988 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3989 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3990 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3991 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3992 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3993 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3994 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3995 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3996 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3997 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3998 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		3999 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4000 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4001 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4002 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4003 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4004 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4005 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4006 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4007 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4008 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4009 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4010 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4011 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4012 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4013 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4014 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4015 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4016 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4017 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4018 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4019 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4020 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4021 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4022 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4023 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4024 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4025 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4026 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4027 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4028 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4029 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4030 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4031 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4032 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4033 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4034 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4035 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4036 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4037 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4038 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4039 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4040 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4041 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4042 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4043 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4044 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4045 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4046 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4047 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4048 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4049 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4050 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4051 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4052 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4053 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4054 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4055 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4056 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4057 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4058 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4059 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4060 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4061 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4062 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4063 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4064 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4065 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4066 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4067 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4068 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4069 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4070 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4071 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4072 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4073 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4074 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4075 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4076 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4077 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4078 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4079 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4080 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4081 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4082 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4083 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4084 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4085 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4086 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4087 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4088 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4089 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4090 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4091 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4092 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4093 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4094 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4095 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4096 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4097 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4098 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4099 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4100 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4101 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4102 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4103 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4104 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4105 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4106 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4107 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4108 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4109 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4110 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4111 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4112 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4113 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4114 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4115 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4116 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4117 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4118 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4119 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4120 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4121 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4122 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4123 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4124 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4125 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4126 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4127 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4128 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4129 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4130 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4131 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4132 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4133 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4134 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4135 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4136 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4137 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4138 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4139 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4140 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4141 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4142 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4143 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4144 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4145 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4146 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4147 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4148 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4149 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4150 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4151 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4152 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4153 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4154 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4155 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4156 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4157 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4158 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4159 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4160 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4161 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4162 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4163 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4164 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4165 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4166 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4167 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4168 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4169 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4170 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4171 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4172 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4173 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4174 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4175 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4176 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4177 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4178 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4179 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4180 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4181 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4182 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4183 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4184 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4185 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4186 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4187 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4188 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4189 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4190 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4191 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4192 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4193 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4194 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4195 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4196 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4197 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4198 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4199 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4200 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4201 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4202 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4203 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4204 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4205 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4206 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4207 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4208 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4209 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4210 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4211 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4212 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4213 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4214 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4215 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4216 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4217 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4218 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4219 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4220 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4221 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4222 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4223 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4224 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4225 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4226 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4227 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4228 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4229 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4230 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4231 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4232 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4233 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4234 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4235 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4236 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4237 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4238 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4239 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4240 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4241 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4242 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4243 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4244 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4245 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4246 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4247 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4248 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4249 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4250 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4251 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4252 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4253 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4254 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4255 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4256 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4257 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4258 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4259 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4260 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4261 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4262 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4263 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4264 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4265 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4266 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4267 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4268 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4269 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4270 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4271 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4272 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4273 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4274 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4275 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4276 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4277 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4278 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4279 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4280 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4281 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4282 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4283 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4284 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4285 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4286 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4287 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4288 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4289 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4290 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4291 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4292 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4293 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4294 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4295 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4296 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4297 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4298 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4299 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4300 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4301 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4302 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4303 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4304 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4305 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4306 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4307 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4308 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4309 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4310 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4311 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4312 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4313 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4314 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4315 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4316 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4317 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4318 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4319 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4320 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4321 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4322 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4323 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4324 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4325 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4326 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4327 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4328 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4329 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4330 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4331 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4332 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4333 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4334 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4335 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4336 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4337 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4338 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4339 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4340 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4341 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4342 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4343 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4344 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4345 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4346 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4347 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4348 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4349 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4350 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4351 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4352 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4353 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4354 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4355 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4356 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4357 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4358 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4359 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4360 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4361 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4362 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4363 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4364 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4365 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4366 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4367 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4368 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4369 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4370 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4371 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4372 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4373 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4374 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4375 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4376 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4377 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4378 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4379 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4380 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4381 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4382 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4383 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4384 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4385 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4386 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4387 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4388 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4389 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4390 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4391 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4392 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4393 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4394 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4395 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4396 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4397 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4398 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4399 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4400 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4401 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4402 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4403 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4404 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4405 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4406 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4407 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4408 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4409 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4410 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4411 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4412 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4413 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4414 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4415 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4416 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4417 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4418 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4419 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4420 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4421 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4422 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4423 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4424 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4425 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4426 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4427 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4428 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4429 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4430 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4431 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4432 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4433 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4434 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4435 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4436 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4437 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4438 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4439 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4440 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4441 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4442 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4443 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4444 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4445 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4446 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4447 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4448 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4449 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4450 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4451 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4452 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4453 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4454 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4455 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4456 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4457 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4458 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4459 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4460 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4461 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4462 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4463 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4464 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4465 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4466 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4467 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4468 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4469 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4470 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4471 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4472 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4473 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4474 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4475 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4476 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4477 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4478 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4479 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4480 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4481 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4482 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4483 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4484 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4485 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4486 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4487 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4488 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4489 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4490 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4491 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4492 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4493 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4494 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4495 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4496 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4497 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4498 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4499 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4500 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4501 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4502 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4503 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4504 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4505 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4506 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4507 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4508 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4509 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4510 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4511 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4512 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4513 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4514 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4515 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4516 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4517 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4518 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4519 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4520 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4521 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4522 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4523 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4524 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4525 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4526 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4527 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4528 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4529 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4530 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4531 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4532 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4533 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4534 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4535 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4536 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4537 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4538 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4539 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4540 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4541 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4542 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4543 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4544 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4545 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4546 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4547 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4548 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4549 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4550 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4551 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4552 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4553 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4554 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4555 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4556 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4557 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4558 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4559 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4560 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4561 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4562 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4563 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4564 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4565 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4566 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4567 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4568 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4569 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4570 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4571 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4572 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4573 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4574 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4575 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4576 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4577 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4578 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4579 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4580 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4581 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4582 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4583 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4584 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4585 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4586 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4587 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4588 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4589 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4590 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4591 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4592 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4593 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4594 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4595 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4596 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4597 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4598 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4599 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4600 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4601 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4602 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4603 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4604 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4605 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4606 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4607 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4608 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4609 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4610 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4611 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4612 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4613 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4614 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4615 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4616 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4617 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4618 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4619 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4620 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4621 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4622 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4623 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4624 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4625 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4626 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4627 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4628 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4629 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4630 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4631 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4632 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4633 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4634 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4635 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4636 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4637 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4638 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4639 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4640 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4641 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4642 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4643 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4644 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4645 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4646 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4647 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4648 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4649 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4650 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4651 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4652 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4653 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4654 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4655 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4656 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4657 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4658 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4659 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4660 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4661 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4662 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4663 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4664 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4665 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4666 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4667 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4668 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4669 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4670 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4671 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4672 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4673 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4674 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4675 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4676 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4677 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4678 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4679 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4680 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4681 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4682 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4683 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4684 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4685 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4686 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4687 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4688 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4689 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4690 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4691 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4692 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4693 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4694 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4695 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4696 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4697 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4698 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4699 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4700 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4701 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4702 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4703 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4704 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4705 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4706 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4707 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4708 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4709 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4710 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4711 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4712 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4713 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4714 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4715 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4716 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4717 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4718 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4719 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4720 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4721 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4722 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4723 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4724 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4725 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4726 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4727 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4728 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4729 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4730 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4731 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4732 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4733 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4734 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4735 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4736 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4737 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4738 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4739 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4740 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4741 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4742 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4743 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4744 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4745 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4746 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4747 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4748 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4749 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4750 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4751 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4752 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4753 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4754 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4755 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4756 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4757 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4758 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4759 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4760 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4761 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4762 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4763 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4764 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4765 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4766 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4767 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4768 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4769 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4770 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4771 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4772 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4773 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4774 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4775 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4776 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4777 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4778 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4779 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4780 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4781 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4782 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4783 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4784 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4785 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4786 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4787 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4788 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4789 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4790 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4791 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4792 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4793 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4794 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4795 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4796 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4797 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4798 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4799 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4800 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4801 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4802 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4803 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4804 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4805 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4806 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4807 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4808 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4809 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4810 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4811 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4812 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4813 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4814 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4815 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4816 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4817 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4818 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4819 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4820 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4821 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4822 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4823 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4824 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4825 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4826 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4827 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4828 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4829 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4830 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4831 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4832 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4833 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4834 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4835 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4836 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4837 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4838 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4839 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4840 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4841 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4842 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4843 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4844 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4845 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4846 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4847 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4848 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4849 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4850 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4851 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4852 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4853 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4854 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4855 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4856 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4857 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4858 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4859 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4860 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4861 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4862 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4863 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4864 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4865 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4866 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4867 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4868 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4869 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4870 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4871 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4872 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4873 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4874 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4875 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4876 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4877 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4878 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4879 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4880 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4881 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4882 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4883 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4884 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4885 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4886 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4887 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4888 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4889 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4890 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4891 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4892 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4893 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4894 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4895 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4896 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4897 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4898 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4899 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4900 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4901 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4902 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4903 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4904 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4905 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4906 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4907 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4908 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4909 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4910 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4911 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4912 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4913 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4914 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4915 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4916 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4917 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4918 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4919 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4920 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4921 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4922 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4923 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4924 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4925 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4926 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4927 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4928 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4929 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4930 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4931 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4932 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4933 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4934 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4935 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4936 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4937 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4938 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4939 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4940 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4941 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4942 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4943 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4944 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4945 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4946 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4947 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4948 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4949 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4950 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4951 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4952 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4953 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4954 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4955 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4956 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4957 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4958 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4959 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4960 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4961 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4962 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4963 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4964 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4965 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4966 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4967 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4968 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4969 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4970 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4971 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4972 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4973 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4974 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4975 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4976 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4977 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4978 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4979 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4980 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4981 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4982 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4983 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4984 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4985 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4986 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4987 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4988 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4989 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4990 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4991 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4992 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4993 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4994 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4995 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4996 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4997 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4998 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		4999 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5000 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5001 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5002 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5003 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5004 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5005 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5006 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5007 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5008 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5009 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5010 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5011 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5012 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5013 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5014 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5015 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5016 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5017 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5018 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5019 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5020 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5021 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5022 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5023 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5024 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5025 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5026 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5027 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5028 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5029 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5030 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5031 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5032 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5033 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5034 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5035 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5036 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5037 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5038 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5039 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5040 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5041 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5042 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5043 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5044 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5045 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5046 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5047 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5048 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5049 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5050 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5051 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5052 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5053 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5054 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5055 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5056 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5057 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5058 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5059 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5060 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5061 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5062 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5063 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5064 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5065 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5066 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5067 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5068 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5069 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5070 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5071 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5072 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5073 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5074 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5075 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5076 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5077 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5078 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5079 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5080 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5081 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5082 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5083 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5084 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5085 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5086 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5087 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5088 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5089 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5090 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5091 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5092 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5093 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5094 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5095 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5096 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5097 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5098 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5099 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5100 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5101 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5102 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5103 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5104 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5105 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5106 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5107 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5108 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5109 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5110 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5111 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5112 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5113 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5114 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5115 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5116 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5117 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5118 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5119 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5120 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5121 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5122 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5123 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5124 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5125 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5126 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5127 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5128 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5129 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5130 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5131 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5132 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5133 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5134 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5135 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5136 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5137 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5138 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5139 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5140 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5141 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5142 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5143 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5144 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5145 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5146 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5147 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5148 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5149 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5150 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5151 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5152 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5153 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5154 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5155 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5156 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5157 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5158 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5159 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5160 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5161 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5162 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5163 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5164 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5165 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5166 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5167 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5168 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5169 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5170 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5171 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5172 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5173 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5174 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5175 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5176 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5177 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5178 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5179 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5180 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5181 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5182 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5183 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5184 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5185 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5186 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5187 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5188 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5189 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5190 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5191 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5192 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5193 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5194 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5195 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5196 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5197 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5198 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5199 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5200 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5201 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5202 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5203 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5204 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5205 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5206 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5207 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5208 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5209 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5210 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5211 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5212 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5213 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5214 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5215 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5216 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5217 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5218 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5219 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5220 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5221 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5222 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5223 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5224 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5225 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5226 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5227 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5228 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5229 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5230 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5231 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5232 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5233 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5234 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5235 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5236 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5237 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5238 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5239 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5240 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5241 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5242 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5243 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5244 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5245 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5246 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5247 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5248 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5249 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5250 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5251 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5252 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5253 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5254 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5255 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5256 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5257 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5258 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5259 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5260 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5261 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5262 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5263 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5264 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5265 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5266 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5267 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5268 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5269 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5270 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5271 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5272 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5273 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5274 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5275 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5276 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5277 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5278 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5279 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5280 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5281 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5282 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5283 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5284 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5285 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5286 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5287 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5288 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5289 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5290 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5291 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5292 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5293 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5294 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5295 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5296 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5297 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5298 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5299 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5300 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5301 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5302 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5303 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5304 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5305 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5306 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5307 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5308 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5309 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5310 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5311 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5312 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5313 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5314 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5315 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5316 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5317 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5318 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5319 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5320 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5321 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5322 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5323 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5324 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5325 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5326 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5327 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5328 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5329 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5330 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5331 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5332 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5333 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5334 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5335 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5336 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5337 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5338 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5339 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5340 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5341 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5342 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5343 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5344 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5345 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5346 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5347 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5348 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5349 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5350 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5351 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5352 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5353 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5354 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5355 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5356 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5357 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5358 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5359 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5360 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5361 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5362 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5363 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5364 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5365 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5366 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5367 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5368 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5369 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5370 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5371 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5372 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5373 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5374 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5375 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5376 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5377 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5378 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5379 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5380 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5381 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5382 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5383 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5384 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5385 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5386 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5387 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5388 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5389 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5390 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5391 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5392 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5393 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5394 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5395 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5396 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5397 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5398 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5399 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5400 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5401 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5402 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5403 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5404 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5405 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5406 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5407 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5408 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5409 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5410 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5411 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5412 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5413 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5414 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5415 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5416 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5417 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5418 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5419 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5420 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5421 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5422 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5423 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5424 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5425 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5426 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5427 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5428 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5429 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5430 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5431 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5432 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5433 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5434 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5435 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5436 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5437 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5438 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5439 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5440 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5441 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5442 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5443 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5444 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5445 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5446 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5447 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5448 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5449 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5450 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5451 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5452 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5453 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5454 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5455 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5456 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5457 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5458 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5459 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5460 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5461 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5462 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5463 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5464 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5465 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5466 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5467 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5468 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5469 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5470 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5471 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5472 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5473 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5474 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5475 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5476 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5477 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5478 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5479 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5480 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5481 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5482 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5483 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5484 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5485 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5486 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5487 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5488 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5489 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5490 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5491 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5492 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5493 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5494 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5495 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5496 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5497 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5498 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5499 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5500 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5501 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5502 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5503 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5504 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5505 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5506 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5507 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5508 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5509 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5510 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5511 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5512 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5513 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5514 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5515 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5516 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5517 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5518 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5519 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5520 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5521 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5522 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5523 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5524 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5525 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5526 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5527 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5528 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5529 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5530 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5531 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5532 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5533 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5534 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5535 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5536 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5537 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5538 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5539 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5540 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5541 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5542 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5543 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5544 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5545 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5546 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5547 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5548 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5549 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5550 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5551 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5552 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5553 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5554 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5555 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5556 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5557 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5558 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5559 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5560 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5561 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5562 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5563 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5564 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5565 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5566 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5567 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5568 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5569 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5570 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5571 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5572 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5573 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5574 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5575 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5576 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5577 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5578 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5579 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5580 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5581 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5582 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5583 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5584 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5585 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5586 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5587 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5588 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5589 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5590 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5591 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5592 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5593 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5594 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5595 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5596 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5597 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5598 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5599 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5600 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5601 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5602 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5603 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5604 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5605 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5606 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5607 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5608 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5609 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5610 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5611 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5612 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5613 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5614 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5615 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5616 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5617 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5618 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5619 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5620 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5621 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5622 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5623 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5624 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5625 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5626 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5627 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5628 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5629 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5630 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5631 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5632 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5633 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5634 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5635 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5636 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5637 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5638 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5639 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5640 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5641 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5642 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5643 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5644 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5645 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5646 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5647 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5648 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5649 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5650 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5651 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5652 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5653 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5654 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5655 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5656 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5657 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5658 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5659 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5660 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5661 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5662 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5663 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5664 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5665 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5666 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5667 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5668 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5669 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5670 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5671 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5672 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5673 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5674 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5675 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5676 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5677 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5678 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5679 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5680 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5681 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5682 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5683 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5684 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5685 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5686 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5687 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5688 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5689 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5690 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5691 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5692 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5693 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5694 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5695 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5696 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5697 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5698 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5699 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5700 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5701 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5702 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5703 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5704 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5705 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5706 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5707 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5708 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5709 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5710 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5711 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5712 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5713 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5714 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5715 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5716 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5717 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5718 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5719 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5720 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5721 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5722 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5723 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5724 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5725 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5726 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5727 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5728 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5729 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5730 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5731 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5732 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5733 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5734 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5735 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5736 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5737 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5738 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5739 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5740 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5741 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5742 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5743 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5744 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5745 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5746 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5747 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5748 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5749 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5750 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5751 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5752 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5753 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5754 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5755 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5756 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5757 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5758 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5759 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5760 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5761 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5762 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5763 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5764 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5765 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5766 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5767 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5768 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5769 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5770 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5771 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5772 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5773 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5774 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5775 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5776 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5777 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5778 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5779 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5780 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5781 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5782 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5783 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5784 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5785 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5786 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5787 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5788 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5789 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5790 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5791 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5792 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5793 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5794 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5795 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5796 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5797 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5798 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5799 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5800 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5801 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5802 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5803 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5804 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5805 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5806 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5807 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5808 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5809 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5810 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5811 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5812 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5813 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5814 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5815 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5816 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5817 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5818 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5819 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5820 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5821 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5822 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5823 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5824 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5825 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5826 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5827 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5828 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5829 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5830 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5831 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5832 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5833 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5834 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5835 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5836 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5837 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5838 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5839 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5840 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5841 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5842 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5843 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5844 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5845 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5846 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5847 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5848 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5849 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5850 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5851 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5852 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5853 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5854 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5855 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5856 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5857 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5858 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5859 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5860 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5861 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5862 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5863 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5864 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5865 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5866 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5867 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5868 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5869 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5870 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5871 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5872 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5873 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5874 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5875 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5876 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5877 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5878 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5879 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5880 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5881 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5882 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5883 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5884 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5885 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5886 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5887 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5888 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5889 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5890 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5891 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5892 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5893 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5894 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5895 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5896 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5897 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5898 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5899 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5900 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5901 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5902 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5903 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5904 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5905 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5906 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5907 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5908 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5909 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5910 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5911 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5912 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5913 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5914 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5915 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5916 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5917 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5918 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5919 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5920 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5921 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5922 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5923 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5924 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5925 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5926 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5927 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5928 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5929 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5930 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5931 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5932 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5933 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5934 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5935 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5936 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5937 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5938 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5939 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5940 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5941 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5942 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5943 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5944 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5945 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5946 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5947 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5948 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5949 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5950 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5951 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5952 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5953 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5954 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5955 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5956 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5957 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5958 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5959 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5960 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5961 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5962 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5963 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5964 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5965 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5966 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5967 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5968 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5969 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5970 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5971 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5972 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5973 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5974 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5975 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5976 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5977 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5978 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5979 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5980 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5981 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5982 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5983 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5984 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5985 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5986 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5987 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5988 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5989 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5990 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5991 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5992 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5993 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5994 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5995 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5996 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5997 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5998 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		5999 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6000 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6001 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6002 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6003 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6004 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6005 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6006 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6007 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6008 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6009 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6010 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6011 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6012 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6013 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6014 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6015 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6016 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6017 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6018 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6019 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6020 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6021 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6022 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6023 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6024 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6025 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6026 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6027 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6028 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6029 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6030 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6031 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6032 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6033 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6034 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6035 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6036 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6037 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6038 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6039 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6040 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6041 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6042 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6043 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6044 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6045 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6046 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6047 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6048 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6049 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6050 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6051 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6052 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6053 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6054 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6055 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6056 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6057 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6058 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6059 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6060 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6061 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6062 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6063 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6064 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6065 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6066 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6067 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6068 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6069 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6070 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6071 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6072 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6073 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6074 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6075 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6076 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6077 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6078 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6079 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6080 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6081 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6082 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6083 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6084 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6085 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6086 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6087 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6088 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6089 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6090 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6091 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6092 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6093 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6094 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6095 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6096 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6097 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6098 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6099 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6100 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6101 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6102 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6103 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6104 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6105 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6106 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6107 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6108 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6109 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6110 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6111 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6112 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6113 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6114 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6115 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6116 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6117 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6118 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6119 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6120 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6121 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6122 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6123 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6124 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6125 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6126 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6127 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6128 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6129 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6130 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6131 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6132 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6133 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6134 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6135 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6136 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6137 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6138 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6139 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6140 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6141 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6142 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6143 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6144 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6145 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6146 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6147 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6148 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6149 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6150 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6151 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6152 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6153 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6154 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6155 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6156 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6157 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6158 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6159 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6160 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6161 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6162 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6163 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6164 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6165 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6166 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6167 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6168 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6169 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6170 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6171 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6172 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6173 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6174 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6175 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6176 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6177 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6178 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6179 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6180 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6181 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6182 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6183 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6184 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6185 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6186 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6187 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6188 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6189 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6190 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6191 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6192 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6193 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6194 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6195 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6196 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6197 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6198 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6199 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6200 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6201 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6202 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6203 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6204 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6205 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6206 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6207 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6208 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6209 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6210 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6211 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6212 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6213 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6214 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6215 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6216 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6217 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6218 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6219 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6220 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6221 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6222 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6223 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6224 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6225 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6226 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6227 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6228 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6229 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6230 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6231 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6232 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6233 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6234 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6235 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6236 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6237 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6238 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6239 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6240 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6241 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6242 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6243 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6244 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6245 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6246 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6247 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6248 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6249 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6250 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6251 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6252 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6253 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6254 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6255 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6256 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6257 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6258 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6259 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6260 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6261 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6262 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6263 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6264 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6265 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6266 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6267 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6268 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6269 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6270 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6271 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6272 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6273 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6274 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6275 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6276 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6277 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6278 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6279 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6280 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6281 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6282 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6283 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6284 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6285 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6286 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6287 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6288 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6289 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6290 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6291 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6292 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6293 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6294 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6295 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6296 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6297 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6298 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6299 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6300 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6301 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6302 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6303 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6304 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6305 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6306 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6307 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6308 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6309 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6310 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6311 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6312 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6313 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6314 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6315 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6316 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6317 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6318 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6319 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6320 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6321 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6322 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6323 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6324 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6325 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6326 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6327 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6328 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6329 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6330 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6331 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6332 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6333 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6334 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6335 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6336 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6337 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6338 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6339 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6340 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6341 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6342 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6343 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6344 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6345 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6346 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6347 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6348 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6349 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6350 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6351 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6352 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6353 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6354 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6355 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6356 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6357 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6358 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6359 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6360 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6361 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6362 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6363 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6364 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6365 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6366 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6367 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6368 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6369 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6370 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6371 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6372 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6373 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6374 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6375 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6376 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6377 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6378 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6379 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6380 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6381 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6382 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6383 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6384 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6385 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6386 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6387 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6388 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6389 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6390 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6391 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6392 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6393 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6394 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6395 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6396 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6397 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6398 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6399 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6400 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6401 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6402 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6403 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6404 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6405 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6406 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6407 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6408 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6409 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6410 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6411 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6412 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6413 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6414 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6415 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6416 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6417 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6418 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6419 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6420 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6421 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6422 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6423 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6424 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6425 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6426 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6427 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6428 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6429 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6430 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6431 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6432 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6433 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6434 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6435 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6436 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6437 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6438 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6439 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6440 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6441 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6442 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6443 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6444 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6445 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6446 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6447 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6448 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6449 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6450 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6451 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6452 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6453 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6454 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6455 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6456 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6457 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6458 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6459 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6460 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6461 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6462 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6463 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6464 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6465 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6466 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6467 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6468 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6469 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6470 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6471 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6472 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6473 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6474 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6475 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6476 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6477 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6478 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6479 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6480 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6481 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6482 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6483 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6484 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6485 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6486 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6487 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6488 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6489 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6490 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6491 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6492 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6493 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6494 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6495 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6496 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6497 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6498 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6499 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6500 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6501 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6502 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6503 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6504 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6505 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6506 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6507 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6508 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6509 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6510 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6511 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6512 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6513 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6514 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6515 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6516 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6517 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6518 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6519 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6520 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6521 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6522 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6523 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6524 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6525 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6526 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6527 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6528 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6529 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6530 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6531 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6532 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6533 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6534 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6535 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6536 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6537 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6538 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6539 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6540 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6541 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6542 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6543 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6544 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6545 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6546 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6547 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6548 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6549 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6550 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6551 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6552 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6553 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6554 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6555 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6556 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6557 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6558 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6559 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6560 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6561 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6562 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6563 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6564 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6565 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6566 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6567 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6568 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6569 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6570 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6571 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6572 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6573 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6574 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6575 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6576 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6577 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6578 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6579 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6580 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6581 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6582 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6583 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6584 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6585 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6586 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6587 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6588 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6589 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6590 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6591 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6592 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6593 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6594 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6595 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6596 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6597 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6598 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6599 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6600 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6601 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6602 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6603 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6604 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6605 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6606 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6607 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6608 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6609 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6610 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6611 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6612 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6613 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6614 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6615 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6616 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6617 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6618 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6619 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6620 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6621 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6622 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6623 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6624 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6625 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6626 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6627 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6628 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6629 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6630 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6631 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6632 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6633 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6634 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6635 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6636 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6637 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6638 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6639 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6640 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6641 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6642 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6643 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6644 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6645 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6646 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6647 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6648 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6649 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6650 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6651 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6652 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6653 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6654 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6655 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6656 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6657 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6658 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6659 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6660 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6661 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6662 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6663 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6664 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6665 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6666 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6667 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6668 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6669 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6670 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6671 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6672 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6673 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6674 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6675 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6676 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6677 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6678 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6679 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6680 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6681 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6682 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6683 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6684 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6685 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6686 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6687 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6688 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6689 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6690 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6691 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6692 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6693 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6694 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6695 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6696 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6697 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6698 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6699 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6700 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6701 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6702 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6703 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6704 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6705 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6706 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6707 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6708 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6709 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6710 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6711 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6712 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6713 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6714 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6715 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6716 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6717 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6718 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6719 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6720 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6721 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6722 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6723 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6724 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6725 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6726 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6727 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6728 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6729 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6730 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6731 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6732 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6733 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6734 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6735 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6736 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6737 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6738 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6739 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6740 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6741 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6742 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6743 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6744 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6745 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6746 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6747 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6748 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6749 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6750 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6751 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6752 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6753 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6754 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6755 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6756 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6757 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6758 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6759 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6760 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6761 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6762 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6763 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6764 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6765 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6766 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6767 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6768 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6769 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6770 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6771 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6772 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6773 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6774 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6775 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6776 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6777 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6778 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6779 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6780 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6781 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6782 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6783 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6784 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6785 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6786 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6787 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6788 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6789 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6790 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6791 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6792 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6793 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6794 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6795 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6796 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6797 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6798 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6799 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6800 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6801 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6802 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6803 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6804 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6805 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6806 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6807 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6808 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6809 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6810 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6811 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6812 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6813 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6814 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6815 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6816 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6817 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6818 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6819 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6820 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6821 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6822 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6823 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6824 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6825 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6826 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6827 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6828 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6829 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6830 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6831 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6832 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6833 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6834 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6835 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6836 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6837 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6838 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6839 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6840 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6841 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6842 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6843 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6844 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6845 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		6846 =>	x"000007BF", -- z: 0 rot: 0 ptr: 1983
		others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;